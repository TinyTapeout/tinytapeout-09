VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_htfab_hybrid
  CLASS BLOCK ;
  FOREIGN tt_um_htfab_hybrid ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.960000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.000000 ;
    ANTENNADIFFAREA 0.478500 ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.000000 ;
    ANTENNADIFFAREA 0.478500 ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.960000 ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.478500 ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.350000 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.350000 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.350000 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.350000 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.350000 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.350000 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.350000 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.350000 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.500000 ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 39.000 5.000 41.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 65.000 5.000 67.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 107.000 5.000 109.000 220.760 ;
    END
  END VAPWR
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 51.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.000 5.000 77.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.000 5.000 119.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.000 5.000 23.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 44.000 5.000 46.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.000 5.000 72.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 112.000 5.000 114.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.000 5.000 18.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 9.000 209.035 29.340 210.465 ;
        RECT 9.000 199.930 10.430 209.035 ;
        RECT 12.430 203.605 25.910 207.035 ;
      LAYER pwell ;
        RECT 12.430 203.355 13.360 203.360 ;
        RECT 12.430 200.575 25.910 203.355 ;
      LAYER nwell ;
        RECT 27.910 199.930 29.340 209.035 ;
        RECT 9.000 198.500 29.340 199.930 ;
        RECT 35.000 208.955 55.340 210.385 ;
        RECT 35.000 193.140 36.430 208.955 ;
      LAYER pwell ;
        RECT 38.430 205.530 51.910 208.310 ;
        RECT 50.980 205.525 51.910 205.530 ;
      LAYER nwell ;
        RECT 38.430 201.850 51.910 205.280 ;
      LAYER pwell ;
        RECT 38.430 198.820 51.910 201.600 ;
        RECT 50.980 198.815 51.910 198.820 ;
      LAYER nwell ;
        RECT 38.430 195.140 51.910 198.570 ;
        RECT 53.910 193.140 55.340 208.955 ;
        RECT 35.000 191.710 55.340 193.140 ;
        RECT 61.000 208.955 81.340 210.385 ;
        RECT 61.000 193.140 62.430 208.955 ;
      LAYER pwell ;
        RECT 64.430 205.530 77.910 208.310 ;
        RECT 76.980 205.525 77.910 205.530 ;
      LAYER nwell ;
        RECT 64.430 201.850 77.910 205.280 ;
      LAYER pwell ;
        RECT 64.430 198.820 77.910 201.600 ;
        RECT 76.980 198.815 77.910 198.820 ;
      LAYER nwell ;
        RECT 64.430 195.140 77.910 198.570 ;
        RECT 79.910 193.140 81.340 208.955 ;
        RECT 103.000 208.955 123.340 210.385 ;
        RECT 103.000 199.850 104.430 208.955 ;
        RECT 106.430 203.525 119.910 206.955 ;
      LAYER pwell ;
        RECT 106.430 203.275 107.360 203.280 ;
        RECT 106.430 200.495 119.910 203.275 ;
      LAYER nwell ;
        RECT 121.910 199.850 123.340 208.955 ;
        RECT 103.000 198.420 123.340 199.850 ;
        RECT 61.000 191.710 81.340 193.140 ;
        RECT 103.000 191.490 123.340 192.920 ;
        RECT 35.000 184.780 55.340 186.210 ;
        RECT 35.000 175.675 36.430 184.780 ;
      LAYER pwell ;
        RECT 38.430 181.355 51.910 184.135 ;
        RECT 50.980 181.350 51.910 181.355 ;
      LAYER nwell ;
        RECT 38.430 177.675 51.910 181.105 ;
        RECT 53.910 175.675 55.340 184.780 ;
        RECT 35.000 174.245 55.340 175.675 ;
        RECT 61.000 184.780 81.340 186.210 ;
        RECT 61.000 175.675 62.430 184.780 ;
      LAYER pwell ;
        RECT 64.430 181.355 77.910 184.135 ;
        RECT 76.980 181.350 77.910 181.355 ;
      LAYER nwell ;
        RECT 64.430 177.675 77.910 181.105 ;
        RECT 79.910 175.675 81.340 184.780 ;
        RECT 61.000 174.245 81.340 175.675 ;
        RECT 103.000 175.675 104.430 191.490 ;
        RECT 106.430 186.060 119.910 189.490 ;
      LAYER pwell ;
        RECT 106.430 185.810 107.360 185.815 ;
        RECT 106.430 183.030 119.910 185.810 ;
      LAYER nwell ;
        RECT 106.430 179.350 119.910 182.780 ;
      LAYER pwell ;
        RECT 106.430 179.100 107.360 179.105 ;
        RECT 106.430 176.320 119.910 179.100 ;
      LAYER nwell ;
        RECT 121.910 175.675 123.340 191.490 ;
        RECT 103.000 174.245 123.340 175.675 ;
        RECT 23.000 149.655 95.355 151.085 ;
        RECT 23.000 130.675 24.430 149.655 ;
        RECT 26.430 132.675 29.860 147.655 ;
      LAYER pwell ;
        RECT 30.110 133.605 32.890 147.655 ;
        RECT 30.105 132.675 32.890 133.605 ;
      LAYER nwell ;
        RECT 33.140 132.675 36.570 147.655 ;
      LAYER pwell ;
        RECT 36.820 133.605 39.600 147.655 ;
        RECT 36.815 132.675 39.600 133.605 ;
      LAYER nwell ;
        RECT 39.850 132.675 43.280 147.655 ;
      LAYER pwell ;
        RECT 43.530 133.605 46.310 147.655 ;
        RECT 43.525 132.675 46.310 133.605 ;
      LAYER nwell ;
        RECT 46.560 132.675 49.990 147.655 ;
      LAYER pwell ;
        RECT 50.240 133.605 53.020 147.655 ;
        RECT 50.235 132.675 53.020 133.605 ;
      LAYER nwell ;
        RECT 53.270 132.675 56.700 147.655 ;
      LAYER pwell ;
        RECT 56.950 133.605 59.730 147.655 ;
        RECT 56.945 132.675 59.730 133.605 ;
      LAYER nwell ;
        RECT 59.980 132.675 63.410 147.655 ;
      LAYER pwell ;
        RECT 63.660 133.605 66.440 147.655 ;
        RECT 63.655 132.675 66.440 133.605 ;
      LAYER nwell ;
        RECT 66.690 132.675 70.120 147.655 ;
      LAYER pwell ;
        RECT 70.370 133.605 73.150 147.655 ;
        RECT 70.365 132.675 73.150 133.605 ;
      LAYER nwell ;
        RECT 73.400 132.675 76.830 147.655 ;
      LAYER pwell ;
        RECT 77.080 133.605 79.860 147.655 ;
        RECT 77.075 132.675 79.860 133.605 ;
      LAYER nwell ;
        RECT 80.110 132.675 83.540 147.655 ;
      LAYER pwell ;
        RECT 83.790 133.605 86.570 147.655 ;
        RECT 83.785 132.675 86.570 133.605 ;
      LAYER nwell ;
        RECT 86.820 132.675 90.250 147.655 ;
      LAYER pwell ;
        RECT 90.500 133.605 93.280 147.655 ;
        RECT 90.495 132.675 93.280 133.605 ;
      LAYER nwell ;
        RECT 93.925 130.675 95.355 149.655 ;
        RECT 23.000 129.245 95.355 130.675 ;
        RECT 29.300 103.140 73.420 104.570 ;
        RECT 29.300 21.430 30.730 103.140 ;
        RECT 32.730 97.710 47.710 101.140 ;
      LAYER pwell ;
        RECT 32.730 97.460 33.660 97.465 ;
        RECT 32.730 94.680 47.710 97.460 ;
      LAYER nwell ;
        RECT 32.730 91.000 47.710 94.430 ;
        RECT 54.705 90.810 69.985 96.420 ;
      LAYER pwell ;
        RECT 32.730 90.750 33.660 90.755 ;
        RECT 32.730 87.970 47.710 90.750 ;
      LAYER nwell ;
        RECT 32.730 84.290 47.710 87.720 ;
      LAYER pwell ;
        RECT 54.705 86.040 69.935 90.560 ;
        RECT 32.730 84.040 33.660 84.045 ;
        RECT 32.730 81.260 47.710 84.040 ;
      LAYER nwell ;
        RECT 32.730 77.580 47.710 81.010 ;
      LAYER pwell ;
        RECT 32.730 77.330 33.660 77.335 ;
        RECT 32.730 74.550 47.710 77.330 ;
      LAYER nwell ;
        RECT 32.730 70.870 47.710 74.300 ;
      LAYER pwell ;
        RECT 32.730 70.620 33.660 70.625 ;
        RECT 32.730 67.840 47.710 70.620 ;
      LAYER nwell ;
        RECT 32.730 64.160 47.710 67.590 ;
      LAYER pwell ;
        RECT 32.730 63.910 33.660 63.915 ;
        RECT 32.730 61.130 47.710 63.910 ;
      LAYER nwell ;
        RECT 32.730 57.450 47.710 60.880 ;
      LAYER pwell ;
        RECT 32.730 57.200 33.660 57.205 ;
        RECT 32.730 54.420 47.710 57.200 ;
      LAYER nwell ;
        RECT 32.730 50.740 47.710 54.170 ;
      LAYER pwell ;
        RECT 32.730 50.490 33.660 50.495 ;
        RECT 32.730 47.710 47.710 50.490 ;
      LAYER nwell ;
        RECT 32.730 44.030 47.710 47.460 ;
      LAYER pwell ;
        RECT 32.730 43.780 33.660 43.785 ;
        RECT 32.730 41.000 47.710 43.780 ;
      LAYER nwell ;
        RECT 54.710 43.775 69.990 49.385 ;
        RECT 32.730 37.320 47.710 40.750 ;
      LAYER pwell ;
        RECT 54.710 39.005 69.940 43.525 ;
      LAYER nwell ;
        RECT 55.350 37.775 67.030 38.755 ;
      LAYER pwell ;
        RECT 32.730 37.070 33.660 37.075 ;
        RECT 32.730 34.290 47.710 37.070 ;
      LAYER nwell ;
        RECT 55.350 27.995 67.010 37.775 ;
        RECT 71.990 21.430 73.420 103.140 ;
        RECT 99.635 74.760 123.005 76.190 ;
        RECT 29.300 20.000 73.420 21.430 ;
        RECT 82.000 34.455 91.720 35.885 ;
        RECT 82.000 21.430 83.430 34.455 ;
        RECT 85.430 26.845 88.290 32.455 ;
      LAYER pwell ;
        RECT 85.430 22.075 88.305 26.600 ;
      LAYER nwell ;
        RECT 90.290 21.430 91.720 34.455 ;
        RECT 82.000 20.000 91.720 21.430 ;
        RECT 99.635 21.430 101.065 74.760 ;
        RECT 105.185 37.775 116.865 38.755 ;
        RECT 105.205 27.995 116.865 37.775 ;
        RECT 121.575 21.430 123.005 74.760 ;
        RECT 99.635 20.000 123.005 21.430 ;
      LAYER li1 ;
        RECT 9.285 210.010 29.055 210.180 ;
        RECT 9.285 198.955 9.455 210.010 ;
        RECT 12.820 206.475 25.520 206.645 ;
        RECT 12.820 204.165 12.990 206.475 ;
        RECT 13.670 206.055 14.170 206.225 ;
        RECT 15.170 206.055 15.670 206.225 ;
        RECT 16.670 206.055 17.170 206.225 ;
        RECT 18.170 206.055 18.670 206.225 ;
        RECT 19.670 206.055 20.170 206.225 ;
        RECT 21.170 206.055 21.670 206.225 ;
        RECT 22.670 206.055 23.170 206.225 ;
        RECT 24.170 206.055 24.670 206.225 ;
        RECT 13.380 204.800 13.550 205.840 ;
        RECT 14.290 204.800 14.460 205.840 ;
        RECT 14.880 204.800 15.050 205.840 ;
        RECT 15.790 204.800 15.960 205.840 ;
        RECT 16.380 204.800 16.550 205.840 ;
        RECT 17.290 204.800 17.460 205.840 ;
        RECT 17.880 204.800 18.050 205.840 ;
        RECT 18.790 204.800 18.960 205.840 ;
        RECT 19.380 204.800 19.550 205.840 ;
        RECT 20.290 204.800 20.460 205.840 ;
        RECT 20.880 204.800 21.050 205.840 ;
        RECT 21.790 204.800 21.960 205.840 ;
        RECT 22.380 204.800 22.550 205.840 ;
        RECT 23.290 204.800 23.460 205.840 ;
        RECT 23.880 204.800 24.050 205.840 ;
        RECT 24.790 204.800 24.960 205.840 ;
        RECT 13.670 204.415 14.170 204.585 ;
        RECT 15.170 204.415 15.670 204.585 ;
        RECT 16.670 204.415 17.170 204.585 ;
        RECT 18.170 204.415 18.670 204.585 ;
        RECT 19.670 204.415 20.170 204.585 ;
        RECT 21.170 204.415 21.670 204.585 ;
        RECT 22.670 204.415 23.170 204.585 ;
        RECT 24.170 204.415 24.670 204.585 ;
        RECT 25.350 204.165 25.520 206.475 ;
        RECT 12.820 203.995 25.520 204.165 ;
        RECT 12.720 202.945 25.670 203.115 ;
        RECT 12.720 200.985 12.890 202.945 ;
        RECT 13.670 202.480 14.170 202.650 ;
        RECT 15.170 202.480 15.670 202.650 ;
        RECT 16.670 202.480 17.170 202.650 ;
        RECT 18.170 202.480 18.670 202.650 ;
        RECT 19.670 202.480 20.170 202.650 ;
        RECT 21.170 202.480 21.670 202.650 ;
        RECT 22.670 202.480 23.170 202.650 ;
        RECT 24.170 202.480 24.670 202.650 ;
        RECT 13.380 201.620 13.550 202.310 ;
        RECT 14.290 201.620 14.460 202.310 ;
        RECT 14.880 201.620 15.050 202.310 ;
        RECT 15.790 201.620 15.960 202.310 ;
        RECT 16.380 201.620 16.550 202.310 ;
        RECT 17.290 201.620 17.460 202.310 ;
        RECT 17.880 201.620 18.050 202.310 ;
        RECT 18.790 201.620 18.960 202.310 ;
        RECT 19.380 201.620 19.550 202.310 ;
        RECT 20.290 201.620 20.460 202.310 ;
        RECT 20.880 201.620 21.050 202.310 ;
        RECT 21.790 201.620 21.960 202.310 ;
        RECT 22.380 201.620 22.550 202.310 ;
        RECT 23.290 201.620 23.460 202.310 ;
        RECT 23.880 201.620 24.050 202.310 ;
        RECT 24.790 201.620 24.960 202.310 ;
        RECT 13.670 201.280 14.170 201.450 ;
        RECT 15.170 201.280 15.670 201.450 ;
        RECT 16.670 201.280 17.170 201.450 ;
        RECT 18.170 201.280 18.670 201.450 ;
        RECT 19.670 201.280 20.170 201.450 ;
        RECT 21.170 201.280 21.670 201.450 ;
        RECT 22.670 201.280 23.170 201.450 ;
        RECT 24.170 201.280 24.670 201.450 ;
        RECT 25.500 200.985 25.670 202.945 ;
        RECT 12.720 200.815 25.670 200.985 ;
        RECT 28.885 198.955 29.055 210.010 ;
        RECT 9.285 198.785 29.055 198.955 ;
        RECT 35.285 209.930 55.055 210.100 ;
        RECT 35.285 192.165 35.455 209.930 ;
        RECT 38.670 207.900 51.620 208.070 ;
        RECT 38.670 205.940 38.840 207.900 ;
        RECT 39.670 207.435 40.170 207.605 ;
        RECT 41.170 207.435 41.670 207.605 ;
        RECT 42.670 207.435 43.170 207.605 ;
        RECT 44.170 207.435 44.670 207.605 ;
        RECT 45.670 207.435 46.170 207.605 ;
        RECT 47.170 207.435 47.670 207.605 ;
        RECT 48.670 207.435 49.170 207.605 ;
        RECT 50.170 207.435 50.670 207.605 ;
        RECT 39.380 206.575 39.550 207.265 ;
        RECT 40.290 206.575 40.460 207.265 ;
        RECT 40.880 206.575 41.050 207.265 ;
        RECT 41.790 206.575 41.960 207.265 ;
        RECT 42.380 206.575 42.550 207.265 ;
        RECT 43.290 206.575 43.460 207.265 ;
        RECT 43.880 206.575 44.050 207.265 ;
        RECT 44.790 206.575 44.960 207.265 ;
        RECT 45.380 206.575 45.550 207.265 ;
        RECT 46.290 206.575 46.460 207.265 ;
        RECT 46.880 206.575 47.050 207.265 ;
        RECT 47.790 206.575 47.960 207.265 ;
        RECT 48.380 206.575 48.550 207.265 ;
        RECT 49.290 206.575 49.460 207.265 ;
        RECT 49.880 206.575 50.050 207.265 ;
        RECT 50.790 206.575 50.960 207.265 ;
        RECT 39.670 206.235 40.170 206.405 ;
        RECT 41.170 206.235 41.670 206.405 ;
        RECT 42.670 206.235 43.170 206.405 ;
        RECT 44.170 206.235 44.670 206.405 ;
        RECT 45.670 206.235 46.170 206.405 ;
        RECT 47.170 206.235 47.670 206.405 ;
        RECT 48.670 206.235 49.170 206.405 ;
        RECT 50.170 206.235 50.670 206.405 ;
        RECT 51.450 205.940 51.620 207.900 ;
        RECT 38.670 205.770 51.620 205.940 ;
        RECT 38.820 204.720 51.520 204.890 ;
        RECT 38.820 202.410 38.990 204.720 ;
        RECT 39.670 204.300 40.170 204.470 ;
        RECT 41.170 204.300 41.670 204.470 ;
        RECT 42.670 204.300 43.170 204.470 ;
        RECT 44.170 204.300 44.670 204.470 ;
        RECT 45.670 204.300 46.170 204.470 ;
        RECT 47.170 204.300 47.670 204.470 ;
        RECT 48.670 204.300 49.170 204.470 ;
        RECT 50.170 204.300 50.670 204.470 ;
        RECT 39.380 203.045 39.550 204.085 ;
        RECT 40.290 203.045 40.460 204.085 ;
        RECT 40.880 203.045 41.050 204.085 ;
        RECT 41.790 203.045 41.960 204.085 ;
        RECT 42.380 203.045 42.550 204.085 ;
        RECT 43.290 203.045 43.460 204.085 ;
        RECT 43.880 203.045 44.050 204.085 ;
        RECT 44.790 203.045 44.960 204.085 ;
        RECT 45.380 203.045 45.550 204.085 ;
        RECT 46.290 203.045 46.460 204.085 ;
        RECT 46.880 203.045 47.050 204.085 ;
        RECT 47.790 203.045 47.960 204.085 ;
        RECT 48.380 203.045 48.550 204.085 ;
        RECT 49.290 203.045 49.460 204.085 ;
        RECT 49.880 203.045 50.050 204.085 ;
        RECT 50.790 203.045 50.960 204.085 ;
        RECT 39.670 202.660 40.170 202.830 ;
        RECT 41.170 202.660 41.670 202.830 ;
        RECT 42.670 202.660 43.170 202.830 ;
        RECT 44.170 202.660 44.670 202.830 ;
        RECT 45.670 202.660 46.170 202.830 ;
        RECT 47.170 202.660 47.670 202.830 ;
        RECT 48.670 202.660 49.170 202.830 ;
        RECT 50.170 202.660 50.670 202.830 ;
        RECT 51.350 202.410 51.520 204.720 ;
        RECT 38.820 202.240 51.520 202.410 ;
        RECT 38.670 201.190 51.620 201.360 ;
        RECT 38.670 199.230 38.840 201.190 ;
        RECT 39.670 200.725 40.170 200.895 ;
        RECT 41.170 200.725 41.670 200.895 ;
        RECT 42.670 200.725 43.170 200.895 ;
        RECT 44.170 200.725 44.670 200.895 ;
        RECT 45.670 200.725 46.170 200.895 ;
        RECT 47.170 200.725 47.670 200.895 ;
        RECT 48.670 200.725 49.170 200.895 ;
        RECT 50.170 200.725 50.670 200.895 ;
        RECT 39.380 199.865 39.550 200.555 ;
        RECT 40.290 199.865 40.460 200.555 ;
        RECT 40.880 199.865 41.050 200.555 ;
        RECT 41.790 199.865 41.960 200.555 ;
        RECT 42.380 199.865 42.550 200.555 ;
        RECT 43.290 199.865 43.460 200.555 ;
        RECT 43.880 199.865 44.050 200.555 ;
        RECT 44.790 199.865 44.960 200.555 ;
        RECT 45.380 199.865 45.550 200.555 ;
        RECT 46.290 199.865 46.460 200.555 ;
        RECT 46.880 199.865 47.050 200.555 ;
        RECT 47.790 199.865 47.960 200.555 ;
        RECT 48.380 199.865 48.550 200.555 ;
        RECT 49.290 199.865 49.460 200.555 ;
        RECT 49.880 199.865 50.050 200.555 ;
        RECT 50.790 199.865 50.960 200.555 ;
        RECT 39.670 199.525 40.170 199.695 ;
        RECT 41.170 199.525 41.670 199.695 ;
        RECT 42.670 199.525 43.170 199.695 ;
        RECT 44.170 199.525 44.670 199.695 ;
        RECT 45.670 199.525 46.170 199.695 ;
        RECT 47.170 199.525 47.670 199.695 ;
        RECT 48.670 199.525 49.170 199.695 ;
        RECT 50.170 199.525 50.670 199.695 ;
        RECT 51.450 199.230 51.620 201.190 ;
        RECT 38.670 199.060 51.620 199.230 ;
        RECT 38.820 198.010 51.520 198.180 ;
        RECT 38.820 195.700 38.990 198.010 ;
        RECT 39.670 197.590 40.170 197.760 ;
        RECT 41.170 197.590 41.670 197.760 ;
        RECT 42.670 197.590 43.170 197.760 ;
        RECT 44.170 197.590 44.670 197.760 ;
        RECT 45.670 197.590 46.170 197.760 ;
        RECT 47.170 197.590 47.670 197.760 ;
        RECT 48.670 197.590 49.170 197.760 ;
        RECT 50.170 197.590 50.670 197.760 ;
        RECT 39.380 196.335 39.550 197.375 ;
        RECT 40.290 196.335 40.460 197.375 ;
        RECT 40.880 196.335 41.050 197.375 ;
        RECT 41.790 196.335 41.960 197.375 ;
        RECT 42.380 196.335 42.550 197.375 ;
        RECT 43.290 196.335 43.460 197.375 ;
        RECT 43.880 196.335 44.050 197.375 ;
        RECT 44.790 196.335 44.960 197.375 ;
        RECT 45.380 196.335 45.550 197.375 ;
        RECT 46.290 196.335 46.460 197.375 ;
        RECT 46.880 196.335 47.050 197.375 ;
        RECT 47.790 196.335 47.960 197.375 ;
        RECT 48.380 196.335 48.550 197.375 ;
        RECT 49.290 196.335 49.460 197.375 ;
        RECT 49.880 196.335 50.050 197.375 ;
        RECT 50.790 196.335 50.960 197.375 ;
        RECT 39.670 195.950 40.170 196.120 ;
        RECT 41.170 195.950 41.670 196.120 ;
        RECT 42.670 195.950 43.170 196.120 ;
        RECT 44.170 195.950 44.670 196.120 ;
        RECT 45.670 195.950 46.170 196.120 ;
        RECT 47.170 195.950 47.670 196.120 ;
        RECT 48.670 195.950 49.170 196.120 ;
        RECT 50.170 195.950 50.670 196.120 ;
        RECT 51.350 195.700 51.520 198.010 ;
        RECT 38.820 195.530 51.520 195.700 ;
        RECT 54.885 192.165 55.055 209.930 ;
        RECT 35.285 191.995 55.055 192.165 ;
        RECT 61.285 209.930 81.055 210.100 ;
        RECT 61.285 192.165 61.455 209.930 ;
        RECT 64.670 207.900 77.620 208.070 ;
        RECT 64.670 205.940 64.840 207.900 ;
        RECT 65.670 207.435 66.170 207.605 ;
        RECT 67.170 207.435 67.670 207.605 ;
        RECT 68.670 207.435 69.170 207.605 ;
        RECT 70.170 207.435 70.670 207.605 ;
        RECT 71.670 207.435 72.170 207.605 ;
        RECT 73.170 207.435 73.670 207.605 ;
        RECT 74.670 207.435 75.170 207.605 ;
        RECT 76.170 207.435 76.670 207.605 ;
        RECT 65.380 206.575 65.550 207.265 ;
        RECT 66.290 206.575 66.460 207.265 ;
        RECT 66.880 206.575 67.050 207.265 ;
        RECT 67.790 206.575 67.960 207.265 ;
        RECT 68.380 206.575 68.550 207.265 ;
        RECT 69.290 206.575 69.460 207.265 ;
        RECT 69.880 206.575 70.050 207.265 ;
        RECT 70.790 206.575 70.960 207.265 ;
        RECT 71.380 206.575 71.550 207.265 ;
        RECT 72.290 206.575 72.460 207.265 ;
        RECT 72.880 206.575 73.050 207.265 ;
        RECT 73.790 206.575 73.960 207.265 ;
        RECT 74.380 206.575 74.550 207.265 ;
        RECT 75.290 206.575 75.460 207.265 ;
        RECT 75.880 206.575 76.050 207.265 ;
        RECT 76.790 206.575 76.960 207.265 ;
        RECT 65.670 206.235 66.170 206.405 ;
        RECT 67.170 206.235 67.670 206.405 ;
        RECT 68.670 206.235 69.170 206.405 ;
        RECT 70.170 206.235 70.670 206.405 ;
        RECT 71.670 206.235 72.170 206.405 ;
        RECT 73.170 206.235 73.670 206.405 ;
        RECT 74.670 206.235 75.170 206.405 ;
        RECT 76.170 206.235 76.670 206.405 ;
        RECT 77.450 205.940 77.620 207.900 ;
        RECT 64.670 205.770 77.620 205.940 ;
        RECT 64.820 204.720 77.520 204.890 ;
        RECT 64.820 202.410 64.990 204.720 ;
        RECT 65.670 204.300 66.170 204.470 ;
        RECT 67.170 204.300 67.670 204.470 ;
        RECT 68.670 204.300 69.170 204.470 ;
        RECT 70.170 204.300 70.670 204.470 ;
        RECT 71.670 204.300 72.170 204.470 ;
        RECT 73.170 204.300 73.670 204.470 ;
        RECT 74.670 204.300 75.170 204.470 ;
        RECT 76.170 204.300 76.670 204.470 ;
        RECT 65.380 203.045 65.550 204.085 ;
        RECT 66.290 203.045 66.460 204.085 ;
        RECT 66.880 203.045 67.050 204.085 ;
        RECT 67.790 203.045 67.960 204.085 ;
        RECT 68.380 203.045 68.550 204.085 ;
        RECT 69.290 203.045 69.460 204.085 ;
        RECT 69.880 203.045 70.050 204.085 ;
        RECT 70.790 203.045 70.960 204.085 ;
        RECT 71.380 203.045 71.550 204.085 ;
        RECT 72.290 203.045 72.460 204.085 ;
        RECT 72.880 203.045 73.050 204.085 ;
        RECT 73.790 203.045 73.960 204.085 ;
        RECT 74.380 203.045 74.550 204.085 ;
        RECT 75.290 203.045 75.460 204.085 ;
        RECT 75.880 203.045 76.050 204.085 ;
        RECT 76.790 203.045 76.960 204.085 ;
        RECT 65.670 202.660 66.170 202.830 ;
        RECT 67.170 202.660 67.670 202.830 ;
        RECT 68.670 202.660 69.170 202.830 ;
        RECT 70.170 202.660 70.670 202.830 ;
        RECT 71.670 202.660 72.170 202.830 ;
        RECT 73.170 202.660 73.670 202.830 ;
        RECT 74.670 202.660 75.170 202.830 ;
        RECT 76.170 202.660 76.670 202.830 ;
        RECT 77.350 202.410 77.520 204.720 ;
        RECT 64.820 202.240 77.520 202.410 ;
        RECT 64.670 201.190 77.620 201.360 ;
        RECT 64.670 199.230 64.840 201.190 ;
        RECT 65.670 200.725 66.170 200.895 ;
        RECT 67.170 200.725 67.670 200.895 ;
        RECT 68.670 200.725 69.170 200.895 ;
        RECT 70.170 200.725 70.670 200.895 ;
        RECT 71.670 200.725 72.170 200.895 ;
        RECT 73.170 200.725 73.670 200.895 ;
        RECT 74.670 200.725 75.170 200.895 ;
        RECT 76.170 200.725 76.670 200.895 ;
        RECT 65.380 199.865 65.550 200.555 ;
        RECT 66.290 199.865 66.460 200.555 ;
        RECT 66.880 199.865 67.050 200.555 ;
        RECT 67.790 199.865 67.960 200.555 ;
        RECT 68.380 199.865 68.550 200.555 ;
        RECT 69.290 199.865 69.460 200.555 ;
        RECT 69.880 199.865 70.050 200.555 ;
        RECT 70.790 199.865 70.960 200.555 ;
        RECT 71.380 199.865 71.550 200.555 ;
        RECT 72.290 199.865 72.460 200.555 ;
        RECT 72.880 199.865 73.050 200.555 ;
        RECT 73.790 199.865 73.960 200.555 ;
        RECT 74.380 199.865 74.550 200.555 ;
        RECT 75.290 199.865 75.460 200.555 ;
        RECT 75.880 199.865 76.050 200.555 ;
        RECT 76.790 199.865 76.960 200.555 ;
        RECT 65.670 199.525 66.170 199.695 ;
        RECT 67.170 199.525 67.670 199.695 ;
        RECT 68.670 199.525 69.170 199.695 ;
        RECT 70.170 199.525 70.670 199.695 ;
        RECT 71.670 199.525 72.170 199.695 ;
        RECT 73.170 199.525 73.670 199.695 ;
        RECT 74.670 199.525 75.170 199.695 ;
        RECT 76.170 199.525 76.670 199.695 ;
        RECT 77.450 199.230 77.620 201.190 ;
        RECT 64.670 199.060 77.620 199.230 ;
        RECT 64.820 198.010 77.520 198.180 ;
        RECT 64.820 195.700 64.990 198.010 ;
        RECT 65.670 197.590 66.170 197.760 ;
        RECT 67.170 197.590 67.670 197.760 ;
        RECT 68.670 197.590 69.170 197.760 ;
        RECT 70.170 197.590 70.670 197.760 ;
        RECT 71.670 197.590 72.170 197.760 ;
        RECT 73.170 197.590 73.670 197.760 ;
        RECT 74.670 197.590 75.170 197.760 ;
        RECT 76.170 197.590 76.670 197.760 ;
        RECT 65.380 196.335 65.550 197.375 ;
        RECT 66.290 196.335 66.460 197.375 ;
        RECT 66.880 196.335 67.050 197.375 ;
        RECT 67.790 196.335 67.960 197.375 ;
        RECT 68.380 196.335 68.550 197.375 ;
        RECT 69.290 196.335 69.460 197.375 ;
        RECT 69.880 196.335 70.050 197.375 ;
        RECT 70.790 196.335 70.960 197.375 ;
        RECT 71.380 196.335 71.550 197.375 ;
        RECT 72.290 196.335 72.460 197.375 ;
        RECT 72.880 196.335 73.050 197.375 ;
        RECT 73.790 196.335 73.960 197.375 ;
        RECT 74.380 196.335 74.550 197.375 ;
        RECT 75.290 196.335 75.460 197.375 ;
        RECT 75.880 196.335 76.050 197.375 ;
        RECT 76.790 196.335 76.960 197.375 ;
        RECT 65.670 195.950 66.170 196.120 ;
        RECT 67.170 195.950 67.670 196.120 ;
        RECT 68.670 195.950 69.170 196.120 ;
        RECT 70.170 195.950 70.670 196.120 ;
        RECT 71.670 195.950 72.170 196.120 ;
        RECT 73.170 195.950 73.670 196.120 ;
        RECT 74.670 195.950 75.170 196.120 ;
        RECT 76.170 195.950 76.670 196.120 ;
        RECT 77.350 195.700 77.520 198.010 ;
        RECT 64.820 195.530 77.520 195.700 ;
        RECT 80.885 192.165 81.055 209.930 ;
        RECT 103.285 209.930 123.055 210.100 ;
        RECT 103.285 198.875 103.455 209.930 ;
        RECT 106.820 206.395 119.520 206.565 ;
        RECT 106.820 204.085 106.990 206.395 ;
        RECT 107.670 205.975 108.170 206.145 ;
        RECT 109.170 205.975 109.670 206.145 ;
        RECT 110.670 205.975 111.170 206.145 ;
        RECT 112.170 205.975 112.670 206.145 ;
        RECT 113.670 205.975 114.170 206.145 ;
        RECT 115.170 205.975 115.670 206.145 ;
        RECT 116.670 205.975 117.170 206.145 ;
        RECT 118.170 205.975 118.670 206.145 ;
        RECT 107.380 204.720 107.550 205.760 ;
        RECT 108.290 204.720 108.460 205.760 ;
        RECT 108.880 204.720 109.050 205.760 ;
        RECT 109.790 204.720 109.960 205.760 ;
        RECT 110.380 204.720 110.550 205.760 ;
        RECT 111.290 204.720 111.460 205.760 ;
        RECT 111.880 204.720 112.050 205.760 ;
        RECT 112.790 204.720 112.960 205.760 ;
        RECT 113.380 204.720 113.550 205.760 ;
        RECT 114.290 204.720 114.460 205.760 ;
        RECT 114.880 204.720 115.050 205.760 ;
        RECT 115.790 204.720 115.960 205.760 ;
        RECT 116.380 204.720 116.550 205.760 ;
        RECT 117.290 204.720 117.460 205.760 ;
        RECT 117.880 204.720 118.050 205.760 ;
        RECT 118.790 204.720 118.960 205.760 ;
        RECT 107.670 204.335 108.170 204.505 ;
        RECT 109.170 204.335 109.670 204.505 ;
        RECT 110.670 204.335 111.170 204.505 ;
        RECT 112.170 204.335 112.670 204.505 ;
        RECT 113.670 204.335 114.170 204.505 ;
        RECT 115.170 204.335 115.670 204.505 ;
        RECT 116.670 204.335 117.170 204.505 ;
        RECT 118.170 204.335 118.670 204.505 ;
        RECT 119.350 204.085 119.520 206.395 ;
        RECT 106.820 203.915 119.520 204.085 ;
        RECT 106.720 202.865 119.670 203.035 ;
        RECT 106.720 200.905 106.890 202.865 ;
        RECT 107.670 202.400 108.170 202.570 ;
        RECT 109.170 202.400 109.670 202.570 ;
        RECT 110.670 202.400 111.170 202.570 ;
        RECT 112.170 202.400 112.670 202.570 ;
        RECT 113.670 202.400 114.170 202.570 ;
        RECT 115.170 202.400 115.670 202.570 ;
        RECT 116.670 202.400 117.170 202.570 ;
        RECT 118.170 202.400 118.670 202.570 ;
        RECT 107.380 201.540 107.550 202.230 ;
        RECT 108.290 201.540 108.460 202.230 ;
        RECT 108.880 201.540 109.050 202.230 ;
        RECT 109.790 201.540 109.960 202.230 ;
        RECT 110.380 201.540 110.550 202.230 ;
        RECT 111.290 201.540 111.460 202.230 ;
        RECT 111.880 201.540 112.050 202.230 ;
        RECT 112.790 201.540 112.960 202.230 ;
        RECT 113.380 201.540 113.550 202.230 ;
        RECT 114.290 201.540 114.460 202.230 ;
        RECT 114.880 201.540 115.050 202.230 ;
        RECT 115.790 201.540 115.960 202.230 ;
        RECT 116.380 201.540 116.550 202.230 ;
        RECT 117.290 201.540 117.460 202.230 ;
        RECT 117.880 201.540 118.050 202.230 ;
        RECT 118.790 201.540 118.960 202.230 ;
        RECT 107.670 201.200 108.170 201.370 ;
        RECT 109.170 201.200 109.670 201.370 ;
        RECT 110.670 201.200 111.170 201.370 ;
        RECT 112.170 201.200 112.670 201.370 ;
        RECT 113.670 201.200 114.170 201.370 ;
        RECT 115.170 201.200 115.670 201.370 ;
        RECT 116.670 201.200 117.170 201.370 ;
        RECT 118.170 201.200 118.670 201.370 ;
        RECT 119.500 200.905 119.670 202.865 ;
        RECT 106.720 200.735 119.670 200.905 ;
        RECT 122.885 198.875 123.055 209.930 ;
        RECT 103.285 198.705 123.055 198.875 ;
        RECT 61.285 191.995 81.055 192.165 ;
        RECT 103.285 192.465 123.055 192.635 ;
        RECT 35.285 185.755 55.055 185.925 ;
        RECT 35.285 174.700 35.455 185.755 ;
        RECT 38.670 183.725 51.620 183.895 ;
        RECT 38.670 181.765 38.840 183.725 ;
        RECT 39.670 183.260 40.170 183.430 ;
        RECT 41.170 183.260 41.670 183.430 ;
        RECT 42.670 183.260 43.170 183.430 ;
        RECT 44.170 183.260 44.670 183.430 ;
        RECT 45.670 183.260 46.170 183.430 ;
        RECT 47.170 183.260 47.670 183.430 ;
        RECT 48.670 183.260 49.170 183.430 ;
        RECT 50.170 183.260 50.670 183.430 ;
        RECT 39.380 182.400 39.550 183.090 ;
        RECT 40.290 182.400 40.460 183.090 ;
        RECT 40.880 182.400 41.050 183.090 ;
        RECT 41.790 182.400 41.960 183.090 ;
        RECT 42.380 182.400 42.550 183.090 ;
        RECT 43.290 182.400 43.460 183.090 ;
        RECT 43.880 182.400 44.050 183.090 ;
        RECT 44.790 182.400 44.960 183.090 ;
        RECT 45.380 182.400 45.550 183.090 ;
        RECT 46.290 182.400 46.460 183.090 ;
        RECT 46.880 182.400 47.050 183.090 ;
        RECT 47.790 182.400 47.960 183.090 ;
        RECT 48.380 182.400 48.550 183.090 ;
        RECT 49.290 182.400 49.460 183.090 ;
        RECT 49.880 182.400 50.050 183.090 ;
        RECT 50.790 182.400 50.960 183.090 ;
        RECT 39.670 182.060 40.170 182.230 ;
        RECT 41.170 182.060 41.670 182.230 ;
        RECT 42.670 182.060 43.170 182.230 ;
        RECT 44.170 182.060 44.670 182.230 ;
        RECT 45.670 182.060 46.170 182.230 ;
        RECT 47.170 182.060 47.670 182.230 ;
        RECT 48.670 182.060 49.170 182.230 ;
        RECT 50.170 182.060 50.670 182.230 ;
        RECT 51.450 181.765 51.620 183.725 ;
        RECT 38.670 181.595 51.620 181.765 ;
        RECT 38.820 180.545 51.520 180.715 ;
        RECT 38.820 178.235 38.990 180.545 ;
        RECT 39.670 180.125 40.170 180.295 ;
        RECT 41.170 180.125 41.670 180.295 ;
        RECT 42.670 180.125 43.170 180.295 ;
        RECT 44.170 180.125 44.670 180.295 ;
        RECT 45.670 180.125 46.170 180.295 ;
        RECT 47.170 180.125 47.670 180.295 ;
        RECT 48.670 180.125 49.170 180.295 ;
        RECT 50.170 180.125 50.670 180.295 ;
        RECT 39.380 178.870 39.550 179.910 ;
        RECT 40.290 178.870 40.460 179.910 ;
        RECT 40.880 178.870 41.050 179.910 ;
        RECT 41.790 178.870 41.960 179.910 ;
        RECT 42.380 178.870 42.550 179.910 ;
        RECT 43.290 178.870 43.460 179.910 ;
        RECT 43.880 178.870 44.050 179.910 ;
        RECT 44.790 178.870 44.960 179.910 ;
        RECT 45.380 178.870 45.550 179.910 ;
        RECT 46.290 178.870 46.460 179.910 ;
        RECT 46.880 178.870 47.050 179.910 ;
        RECT 47.790 178.870 47.960 179.910 ;
        RECT 48.380 178.870 48.550 179.910 ;
        RECT 49.290 178.870 49.460 179.910 ;
        RECT 49.880 178.870 50.050 179.910 ;
        RECT 50.790 178.870 50.960 179.910 ;
        RECT 39.670 178.485 40.170 178.655 ;
        RECT 41.170 178.485 41.670 178.655 ;
        RECT 42.670 178.485 43.170 178.655 ;
        RECT 44.170 178.485 44.670 178.655 ;
        RECT 45.670 178.485 46.170 178.655 ;
        RECT 47.170 178.485 47.670 178.655 ;
        RECT 48.670 178.485 49.170 178.655 ;
        RECT 50.170 178.485 50.670 178.655 ;
        RECT 51.350 178.235 51.520 180.545 ;
        RECT 38.820 178.065 51.520 178.235 ;
        RECT 54.885 174.700 55.055 185.755 ;
        RECT 35.285 174.530 55.055 174.700 ;
        RECT 61.285 185.755 81.055 185.925 ;
        RECT 61.285 174.700 61.455 185.755 ;
        RECT 64.670 183.725 77.620 183.895 ;
        RECT 64.670 181.765 64.840 183.725 ;
        RECT 65.670 183.260 66.170 183.430 ;
        RECT 67.170 183.260 67.670 183.430 ;
        RECT 68.670 183.260 69.170 183.430 ;
        RECT 70.170 183.260 70.670 183.430 ;
        RECT 71.670 183.260 72.170 183.430 ;
        RECT 73.170 183.260 73.670 183.430 ;
        RECT 74.670 183.260 75.170 183.430 ;
        RECT 76.170 183.260 76.670 183.430 ;
        RECT 65.380 182.400 65.550 183.090 ;
        RECT 66.290 182.400 66.460 183.090 ;
        RECT 66.880 182.400 67.050 183.090 ;
        RECT 67.790 182.400 67.960 183.090 ;
        RECT 68.380 182.400 68.550 183.090 ;
        RECT 69.290 182.400 69.460 183.090 ;
        RECT 69.880 182.400 70.050 183.090 ;
        RECT 70.790 182.400 70.960 183.090 ;
        RECT 71.380 182.400 71.550 183.090 ;
        RECT 72.290 182.400 72.460 183.090 ;
        RECT 72.880 182.400 73.050 183.090 ;
        RECT 73.790 182.400 73.960 183.090 ;
        RECT 74.380 182.400 74.550 183.090 ;
        RECT 75.290 182.400 75.460 183.090 ;
        RECT 75.880 182.400 76.050 183.090 ;
        RECT 76.790 182.400 76.960 183.090 ;
        RECT 65.670 182.060 66.170 182.230 ;
        RECT 67.170 182.060 67.670 182.230 ;
        RECT 68.670 182.060 69.170 182.230 ;
        RECT 70.170 182.060 70.670 182.230 ;
        RECT 71.670 182.060 72.170 182.230 ;
        RECT 73.170 182.060 73.670 182.230 ;
        RECT 74.670 182.060 75.170 182.230 ;
        RECT 76.170 182.060 76.670 182.230 ;
        RECT 77.450 181.765 77.620 183.725 ;
        RECT 64.670 181.595 77.620 181.765 ;
        RECT 64.820 180.545 77.520 180.715 ;
        RECT 64.820 178.235 64.990 180.545 ;
        RECT 65.670 180.125 66.170 180.295 ;
        RECT 67.170 180.125 67.670 180.295 ;
        RECT 68.670 180.125 69.170 180.295 ;
        RECT 70.170 180.125 70.670 180.295 ;
        RECT 71.670 180.125 72.170 180.295 ;
        RECT 73.170 180.125 73.670 180.295 ;
        RECT 74.670 180.125 75.170 180.295 ;
        RECT 76.170 180.125 76.670 180.295 ;
        RECT 65.380 178.870 65.550 179.910 ;
        RECT 66.290 178.870 66.460 179.910 ;
        RECT 66.880 178.870 67.050 179.910 ;
        RECT 67.790 178.870 67.960 179.910 ;
        RECT 68.380 178.870 68.550 179.910 ;
        RECT 69.290 178.870 69.460 179.910 ;
        RECT 69.880 178.870 70.050 179.910 ;
        RECT 70.790 178.870 70.960 179.910 ;
        RECT 71.380 178.870 71.550 179.910 ;
        RECT 72.290 178.870 72.460 179.910 ;
        RECT 72.880 178.870 73.050 179.910 ;
        RECT 73.790 178.870 73.960 179.910 ;
        RECT 74.380 178.870 74.550 179.910 ;
        RECT 75.290 178.870 75.460 179.910 ;
        RECT 75.880 178.870 76.050 179.910 ;
        RECT 76.790 178.870 76.960 179.910 ;
        RECT 65.670 178.485 66.170 178.655 ;
        RECT 67.170 178.485 67.670 178.655 ;
        RECT 68.670 178.485 69.170 178.655 ;
        RECT 70.170 178.485 70.670 178.655 ;
        RECT 71.670 178.485 72.170 178.655 ;
        RECT 73.170 178.485 73.670 178.655 ;
        RECT 74.670 178.485 75.170 178.655 ;
        RECT 76.170 178.485 76.670 178.655 ;
        RECT 77.350 178.235 77.520 180.545 ;
        RECT 64.820 178.065 77.520 178.235 ;
        RECT 80.885 174.700 81.055 185.755 ;
        RECT 61.285 174.530 81.055 174.700 ;
        RECT 103.285 174.700 103.455 192.465 ;
        RECT 106.820 188.930 119.520 189.100 ;
        RECT 106.820 186.620 106.990 188.930 ;
        RECT 107.670 188.510 108.170 188.680 ;
        RECT 109.170 188.510 109.670 188.680 ;
        RECT 110.670 188.510 111.170 188.680 ;
        RECT 112.170 188.510 112.670 188.680 ;
        RECT 113.670 188.510 114.170 188.680 ;
        RECT 115.170 188.510 115.670 188.680 ;
        RECT 116.670 188.510 117.170 188.680 ;
        RECT 118.170 188.510 118.670 188.680 ;
        RECT 107.380 187.255 107.550 188.295 ;
        RECT 108.290 187.255 108.460 188.295 ;
        RECT 108.880 187.255 109.050 188.295 ;
        RECT 109.790 187.255 109.960 188.295 ;
        RECT 110.380 187.255 110.550 188.295 ;
        RECT 111.290 187.255 111.460 188.295 ;
        RECT 111.880 187.255 112.050 188.295 ;
        RECT 112.790 187.255 112.960 188.295 ;
        RECT 113.380 187.255 113.550 188.295 ;
        RECT 114.290 187.255 114.460 188.295 ;
        RECT 114.880 187.255 115.050 188.295 ;
        RECT 115.790 187.255 115.960 188.295 ;
        RECT 116.380 187.255 116.550 188.295 ;
        RECT 117.290 187.255 117.460 188.295 ;
        RECT 117.880 187.255 118.050 188.295 ;
        RECT 118.790 187.255 118.960 188.295 ;
        RECT 107.670 186.870 108.170 187.040 ;
        RECT 109.170 186.870 109.670 187.040 ;
        RECT 110.670 186.870 111.170 187.040 ;
        RECT 112.170 186.870 112.670 187.040 ;
        RECT 113.670 186.870 114.170 187.040 ;
        RECT 115.170 186.870 115.670 187.040 ;
        RECT 116.670 186.870 117.170 187.040 ;
        RECT 118.170 186.870 118.670 187.040 ;
        RECT 119.350 186.620 119.520 188.930 ;
        RECT 106.820 186.450 119.520 186.620 ;
        RECT 106.720 185.400 119.670 185.570 ;
        RECT 106.720 183.440 106.890 185.400 ;
        RECT 107.670 184.935 108.170 185.105 ;
        RECT 109.170 184.935 109.670 185.105 ;
        RECT 110.670 184.935 111.170 185.105 ;
        RECT 112.170 184.935 112.670 185.105 ;
        RECT 113.670 184.935 114.170 185.105 ;
        RECT 115.170 184.935 115.670 185.105 ;
        RECT 116.670 184.935 117.170 185.105 ;
        RECT 118.170 184.935 118.670 185.105 ;
        RECT 107.380 184.075 107.550 184.765 ;
        RECT 108.290 184.075 108.460 184.765 ;
        RECT 108.880 184.075 109.050 184.765 ;
        RECT 109.790 184.075 109.960 184.765 ;
        RECT 110.380 184.075 110.550 184.765 ;
        RECT 111.290 184.075 111.460 184.765 ;
        RECT 111.880 184.075 112.050 184.765 ;
        RECT 112.790 184.075 112.960 184.765 ;
        RECT 113.380 184.075 113.550 184.765 ;
        RECT 114.290 184.075 114.460 184.765 ;
        RECT 114.880 184.075 115.050 184.765 ;
        RECT 115.790 184.075 115.960 184.765 ;
        RECT 116.380 184.075 116.550 184.765 ;
        RECT 117.290 184.075 117.460 184.765 ;
        RECT 117.880 184.075 118.050 184.765 ;
        RECT 118.790 184.075 118.960 184.765 ;
        RECT 107.670 183.735 108.170 183.905 ;
        RECT 109.170 183.735 109.670 183.905 ;
        RECT 110.670 183.735 111.170 183.905 ;
        RECT 112.170 183.735 112.670 183.905 ;
        RECT 113.670 183.735 114.170 183.905 ;
        RECT 115.170 183.735 115.670 183.905 ;
        RECT 116.670 183.735 117.170 183.905 ;
        RECT 118.170 183.735 118.670 183.905 ;
        RECT 119.500 183.440 119.670 185.400 ;
        RECT 106.720 183.270 119.670 183.440 ;
        RECT 106.820 182.220 119.520 182.390 ;
        RECT 106.820 179.910 106.990 182.220 ;
        RECT 107.670 181.800 108.170 181.970 ;
        RECT 109.170 181.800 109.670 181.970 ;
        RECT 110.670 181.800 111.170 181.970 ;
        RECT 112.170 181.800 112.670 181.970 ;
        RECT 113.670 181.800 114.170 181.970 ;
        RECT 115.170 181.800 115.670 181.970 ;
        RECT 116.670 181.800 117.170 181.970 ;
        RECT 118.170 181.800 118.670 181.970 ;
        RECT 107.380 180.545 107.550 181.585 ;
        RECT 108.290 180.545 108.460 181.585 ;
        RECT 108.880 180.545 109.050 181.585 ;
        RECT 109.790 180.545 109.960 181.585 ;
        RECT 110.380 180.545 110.550 181.585 ;
        RECT 111.290 180.545 111.460 181.585 ;
        RECT 111.880 180.545 112.050 181.585 ;
        RECT 112.790 180.545 112.960 181.585 ;
        RECT 113.380 180.545 113.550 181.585 ;
        RECT 114.290 180.545 114.460 181.585 ;
        RECT 114.880 180.545 115.050 181.585 ;
        RECT 115.790 180.545 115.960 181.585 ;
        RECT 116.380 180.545 116.550 181.585 ;
        RECT 117.290 180.545 117.460 181.585 ;
        RECT 117.880 180.545 118.050 181.585 ;
        RECT 118.790 180.545 118.960 181.585 ;
        RECT 107.670 180.160 108.170 180.330 ;
        RECT 109.170 180.160 109.670 180.330 ;
        RECT 110.670 180.160 111.170 180.330 ;
        RECT 112.170 180.160 112.670 180.330 ;
        RECT 113.670 180.160 114.170 180.330 ;
        RECT 115.170 180.160 115.670 180.330 ;
        RECT 116.670 180.160 117.170 180.330 ;
        RECT 118.170 180.160 118.670 180.330 ;
        RECT 119.350 179.910 119.520 182.220 ;
        RECT 106.820 179.740 119.520 179.910 ;
        RECT 106.720 178.690 119.670 178.860 ;
        RECT 106.720 176.730 106.890 178.690 ;
        RECT 107.670 178.225 108.170 178.395 ;
        RECT 109.170 178.225 109.670 178.395 ;
        RECT 110.670 178.225 111.170 178.395 ;
        RECT 112.170 178.225 112.670 178.395 ;
        RECT 113.670 178.225 114.170 178.395 ;
        RECT 115.170 178.225 115.670 178.395 ;
        RECT 116.670 178.225 117.170 178.395 ;
        RECT 118.170 178.225 118.670 178.395 ;
        RECT 107.380 177.365 107.550 178.055 ;
        RECT 108.290 177.365 108.460 178.055 ;
        RECT 108.880 177.365 109.050 178.055 ;
        RECT 109.790 177.365 109.960 178.055 ;
        RECT 110.380 177.365 110.550 178.055 ;
        RECT 111.290 177.365 111.460 178.055 ;
        RECT 111.880 177.365 112.050 178.055 ;
        RECT 112.790 177.365 112.960 178.055 ;
        RECT 113.380 177.365 113.550 178.055 ;
        RECT 114.290 177.365 114.460 178.055 ;
        RECT 114.880 177.365 115.050 178.055 ;
        RECT 115.790 177.365 115.960 178.055 ;
        RECT 116.380 177.365 116.550 178.055 ;
        RECT 117.290 177.365 117.460 178.055 ;
        RECT 117.880 177.365 118.050 178.055 ;
        RECT 118.790 177.365 118.960 178.055 ;
        RECT 107.670 177.025 108.170 177.195 ;
        RECT 109.170 177.025 109.670 177.195 ;
        RECT 110.670 177.025 111.170 177.195 ;
        RECT 112.170 177.025 112.670 177.195 ;
        RECT 113.670 177.025 114.170 177.195 ;
        RECT 115.170 177.025 115.670 177.195 ;
        RECT 116.670 177.025 117.170 177.195 ;
        RECT 118.170 177.025 118.670 177.195 ;
        RECT 119.500 176.730 119.670 178.690 ;
        RECT 106.720 176.560 119.670 176.730 ;
        RECT 122.885 174.700 123.055 192.465 ;
        RECT 103.285 174.530 123.055 174.700 ;
        RECT 23.285 150.630 95.070 150.800 ;
        RECT 23.285 129.700 23.455 150.630 ;
        RECT 26.820 147.095 29.470 147.265 ;
        RECT 26.820 133.235 26.990 147.095 ;
        RECT 27.625 146.535 28.665 146.705 ;
        RECT 27.240 145.915 27.410 146.415 ;
        RECT 28.880 145.915 29.050 146.415 ;
        RECT 27.625 145.625 28.665 145.795 ;
        RECT 27.625 145.035 28.665 145.205 ;
        RECT 27.240 144.415 27.410 144.915 ;
        RECT 28.880 144.415 29.050 144.915 ;
        RECT 27.625 144.125 28.665 144.295 ;
        RECT 27.625 143.535 28.665 143.705 ;
        RECT 27.240 142.915 27.410 143.415 ;
        RECT 28.880 142.915 29.050 143.415 ;
        RECT 27.625 142.625 28.665 142.795 ;
        RECT 27.625 142.035 28.665 142.205 ;
        RECT 27.240 141.415 27.410 141.915 ;
        RECT 28.880 141.415 29.050 141.915 ;
        RECT 27.625 141.125 28.665 141.295 ;
        RECT 27.625 140.535 28.665 140.705 ;
        RECT 27.240 139.915 27.410 140.415 ;
        RECT 28.880 139.915 29.050 140.415 ;
        RECT 27.625 139.625 28.665 139.795 ;
        RECT 27.625 139.035 28.665 139.205 ;
        RECT 27.240 138.415 27.410 138.915 ;
        RECT 28.880 138.415 29.050 138.915 ;
        RECT 27.625 138.125 28.665 138.295 ;
        RECT 27.625 137.535 28.665 137.705 ;
        RECT 27.240 136.915 27.410 137.415 ;
        RECT 28.880 136.915 29.050 137.415 ;
        RECT 27.625 136.625 28.665 136.795 ;
        RECT 27.625 136.035 28.665 136.205 ;
        RECT 27.240 135.415 27.410 135.915 ;
        RECT 28.880 135.415 29.050 135.915 ;
        RECT 27.625 135.125 28.665 135.295 ;
        RECT 27.625 134.535 28.665 134.705 ;
        RECT 27.240 133.915 27.410 134.415 ;
        RECT 28.880 133.915 29.050 134.415 ;
        RECT 27.625 133.625 28.665 133.795 ;
        RECT 29.300 133.235 29.470 147.095 ;
        RECT 26.820 133.065 29.470 133.235 ;
        RECT 30.350 147.245 32.650 147.415 ;
        RECT 30.350 133.135 30.520 147.245 ;
        RECT 31.155 146.535 31.845 146.705 ;
        RECT 30.815 145.915 30.985 146.415 ;
        RECT 32.015 145.915 32.185 146.415 ;
        RECT 31.155 145.625 31.845 145.795 ;
        RECT 31.155 145.035 31.845 145.205 ;
        RECT 30.815 144.415 30.985 144.915 ;
        RECT 32.015 144.415 32.185 144.915 ;
        RECT 31.155 144.125 31.845 144.295 ;
        RECT 31.155 143.535 31.845 143.705 ;
        RECT 30.815 142.915 30.985 143.415 ;
        RECT 32.015 142.915 32.185 143.415 ;
        RECT 31.155 142.625 31.845 142.795 ;
        RECT 31.155 142.035 31.845 142.205 ;
        RECT 30.815 141.415 30.985 141.915 ;
        RECT 32.015 141.415 32.185 141.915 ;
        RECT 31.155 141.125 31.845 141.295 ;
        RECT 31.155 140.535 31.845 140.705 ;
        RECT 30.815 139.915 30.985 140.415 ;
        RECT 32.015 139.915 32.185 140.415 ;
        RECT 31.155 139.625 31.845 139.795 ;
        RECT 31.155 139.035 31.845 139.205 ;
        RECT 30.815 138.415 30.985 138.915 ;
        RECT 32.015 138.415 32.185 138.915 ;
        RECT 31.155 138.125 31.845 138.295 ;
        RECT 31.155 137.535 31.845 137.705 ;
        RECT 30.815 136.915 30.985 137.415 ;
        RECT 32.015 136.915 32.185 137.415 ;
        RECT 31.155 136.625 31.845 136.795 ;
        RECT 31.155 136.035 31.845 136.205 ;
        RECT 30.815 135.415 30.985 135.915 ;
        RECT 32.015 135.415 32.185 135.915 ;
        RECT 31.155 135.125 31.845 135.295 ;
        RECT 31.155 134.535 31.845 134.705 ;
        RECT 30.815 133.915 30.985 134.415 ;
        RECT 32.015 133.915 32.185 134.415 ;
        RECT 31.155 133.625 31.845 133.795 ;
        RECT 32.480 133.135 32.650 147.245 ;
        RECT 30.350 132.965 32.650 133.135 ;
        RECT 33.530 147.095 36.180 147.265 ;
        RECT 33.530 133.235 33.700 147.095 ;
        RECT 34.335 146.535 35.375 146.705 ;
        RECT 33.950 145.915 34.120 146.415 ;
        RECT 35.590 145.915 35.760 146.415 ;
        RECT 34.335 145.625 35.375 145.795 ;
        RECT 34.335 145.035 35.375 145.205 ;
        RECT 33.950 144.415 34.120 144.915 ;
        RECT 35.590 144.415 35.760 144.915 ;
        RECT 34.335 144.125 35.375 144.295 ;
        RECT 34.335 143.535 35.375 143.705 ;
        RECT 33.950 142.915 34.120 143.415 ;
        RECT 35.590 142.915 35.760 143.415 ;
        RECT 34.335 142.625 35.375 142.795 ;
        RECT 34.335 142.035 35.375 142.205 ;
        RECT 33.950 141.415 34.120 141.915 ;
        RECT 35.590 141.415 35.760 141.915 ;
        RECT 34.335 141.125 35.375 141.295 ;
        RECT 34.335 140.535 35.375 140.705 ;
        RECT 33.950 139.915 34.120 140.415 ;
        RECT 35.590 139.915 35.760 140.415 ;
        RECT 34.335 139.625 35.375 139.795 ;
        RECT 34.335 139.035 35.375 139.205 ;
        RECT 33.950 138.415 34.120 138.915 ;
        RECT 35.590 138.415 35.760 138.915 ;
        RECT 34.335 138.125 35.375 138.295 ;
        RECT 34.335 137.535 35.375 137.705 ;
        RECT 33.950 136.915 34.120 137.415 ;
        RECT 35.590 136.915 35.760 137.415 ;
        RECT 34.335 136.625 35.375 136.795 ;
        RECT 34.335 136.035 35.375 136.205 ;
        RECT 33.950 135.415 34.120 135.915 ;
        RECT 35.590 135.415 35.760 135.915 ;
        RECT 34.335 135.125 35.375 135.295 ;
        RECT 34.335 134.535 35.375 134.705 ;
        RECT 33.950 133.915 34.120 134.415 ;
        RECT 35.590 133.915 35.760 134.415 ;
        RECT 34.335 133.625 35.375 133.795 ;
        RECT 36.010 133.235 36.180 147.095 ;
        RECT 33.530 133.065 36.180 133.235 ;
        RECT 37.060 147.245 39.360 147.415 ;
        RECT 37.060 133.135 37.230 147.245 ;
        RECT 37.865 146.535 38.555 146.705 ;
        RECT 37.525 145.915 37.695 146.415 ;
        RECT 38.725 145.915 38.895 146.415 ;
        RECT 37.865 145.625 38.555 145.795 ;
        RECT 37.865 145.035 38.555 145.205 ;
        RECT 37.525 144.415 37.695 144.915 ;
        RECT 38.725 144.415 38.895 144.915 ;
        RECT 37.865 144.125 38.555 144.295 ;
        RECT 37.865 143.535 38.555 143.705 ;
        RECT 37.525 142.915 37.695 143.415 ;
        RECT 38.725 142.915 38.895 143.415 ;
        RECT 37.865 142.625 38.555 142.795 ;
        RECT 37.865 142.035 38.555 142.205 ;
        RECT 37.525 141.415 37.695 141.915 ;
        RECT 38.725 141.415 38.895 141.915 ;
        RECT 37.865 141.125 38.555 141.295 ;
        RECT 37.865 140.535 38.555 140.705 ;
        RECT 37.525 139.915 37.695 140.415 ;
        RECT 38.725 139.915 38.895 140.415 ;
        RECT 37.865 139.625 38.555 139.795 ;
        RECT 37.865 139.035 38.555 139.205 ;
        RECT 37.525 138.415 37.695 138.915 ;
        RECT 38.725 138.415 38.895 138.915 ;
        RECT 37.865 138.125 38.555 138.295 ;
        RECT 37.865 137.535 38.555 137.705 ;
        RECT 37.525 136.915 37.695 137.415 ;
        RECT 38.725 136.915 38.895 137.415 ;
        RECT 37.865 136.625 38.555 136.795 ;
        RECT 37.865 136.035 38.555 136.205 ;
        RECT 37.525 135.415 37.695 135.915 ;
        RECT 38.725 135.415 38.895 135.915 ;
        RECT 37.865 135.125 38.555 135.295 ;
        RECT 37.865 134.535 38.555 134.705 ;
        RECT 37.525 133.915 37.695 134.415 ;
        RECT 38.725 133.915 38.895 134.415 ;
        RECT 37.865 133.625 38.555 133.795 ;
        RECT 39.190 133.135 39.360 147.245 ;
        RECT 37.060 132.965 39.360 133.135 ;
        RECT 40.240 147.095 42.890 147.265 ;
        RECT 40.240 133.235 40.410 147.095 ;
        RECT 41.045 146.535 42.085 146.705 ;
        RECT 40.660 145.915 40.830 146.415 ;
        RECT 42.300 145.915 42.470 146.415 ;
        RECT 41.045 145.625 42.085 145.795 ;
        RECT 41.045 145.035 42.085 145.205 ;
        RECT 40.660 144.415 40.830 144.915 ;
        RECT 42.300 144.415 42.470 144.915 ;
        RECT 41.045 144.125 42.085 144.295 ;
        RECT 41.045 143.535 42.085 143.705 ;
        RECT 40.660 142.915 40.830 143.415 ;
        RECT 42.300 142.915 42.470 143.415 ;
        RECT 41.045 142.625 42.085 142.795 ;
        RECT 41.045 142.035 42.085 142.205 ;
        RECT 40.660 141.415 40.830 141.915 ;
        RECT 42.300 141.415 42.470 141.915 ;
        RECT 41.045 141.125 42.085 141.295 ;
        RECT 41.045 140.535 42.085 140.705 ;
        RECT 40.660 139.915 40.830 140.415 ;
        RECT 42.300 139.915 42.470 140.415 ;
        RECT 41.045 139.625 42.085 139.795 ;
        RECT 41.045 139.035 42.085 139.205 ;
        RECT 40.660 138.415 40.830 138.915 ;
        RECT 42.300 138.415 42.470 138.915 ;
        RECT 41.045 138.125 42.085 138.295 ;
        RECT 41.045 137.535 42.085 137.705 ;
        RECT 40.660 136.915 40.830 137.415 ;
        RECT 42.300 136.915 42.470 137.415 ;
        RECT 41.045 136.625 42.085 136.795 ;
        RECT 41.045 136.035 42.085 136.205 ;
        RECT 40.660 135.415 40.830 135.915 ;
        RECT 42.300 135.415 42.470 135.915 ;
        RECT 41.045 135.125 42.085 135.295 ;
        RECT 41.045 134.535 42.085 134.705 ;
        RECT 40.660 133.915 40.830 134.415 ;
        RECT 42.300 133.915 42.470 134.415 ;
        RECT 41.045 133.625 42.085 133.795 ;
        RECT 42.720 133.235 42.890 147.095 ;
        RECT 40.240 133.065 42.890 133.235 ;
        RECT 43.770 147.245 46.070 147.415 ;
        RECT 43.770 133.135 43.940 147.245 ;
        RECT 44.575 146.535 45.265 146.705 ;
        RECT 44.235 145.915 44.405 146.415 ;
        RECT 45.435 145.915 45.605 146.415 ;
        RECT 44.575 145.625 45.265 145.795 ;
        RECT 44.575 145.035 45.265 145.205 ;
        RECT 44.235 144.415 44.405 144.915 ;
        RECT 45.435 144.415 45.605 144.915 ;
        RECT 44.575 144.125 45.265 144.295 ;
        RECT 44.575 143.535 45.265 143.705 ;
        RECT 44.235 142.915 44.405 143.415 ;
        RECT 45.435 142.915 45.605 143.415 ;
        RECT 44.575 142.625 45.265 142.795 ;
        RECT 44.575 142.035 45.265 142.205 ;
        RECT 44.235 141.415 44.405 141.915 ;
        RECT 45.435 141.415 45.605 141.915 ;
        RECT 44.575 141.125 45.265 141.295 ;
        RECT 44.575 140.535 45.265 140.705 ;
        RECT 44.235 139.915 44.405 140.415 ;
        RECT 45.435 139.915 45.605 140.415 ;
        RECT 44.575 139.625 45.265 139.795 ;
        RECT 44.575 139.035 45.265 139.205 ;
        RECT 44.235 138.415 44.405 138.915 ;
        RECT 45.435 138.415 45.605 138.915 ;
        RECT 44.575 138.125 45.265 138.295 ;
        RECT 44.575 137.535 45.265 137.705 ;
        RECT 44.235 136.915 44.405 137.415 ;
        RECT 45.435 136.915 45.605 137.415 ;
        RECT 44.575 136.625 45.265 136.795 ;
        RECT 44.575 136.035 45.265 136.205 ;
        RECT 44.235 135.415 44.405 135.915 ;
        RECT 45.435 135.415 45.605 135.915 ;
        RECT 44.575 135.125 45.265 135.295 ;
        RECT 44.575 134.535 45.265 134.705 ;
        RECT 44.235 133.915 44.405 134.415 ;
        RECT 45.435 133.915 45.605 134.415 ;
        RECT 44.575 133.625 45.265 133.795 ;
        RECT 45.900 133.135 46.070 147.245 ;
        RECT 43.770 132.965 46.070 133.135 ;
        RECT 46.950 147.095 49.600 147.265 ;
        RECT 46.950 133.235 47.120 147.095 ;
        RECT 47.755 146.535 48.795 146.705 ;
        RECT 47.370 145.915 47.540 146.415 ;
        RECT 49.010 145.915 49.180 146.415 ;
        RECT 47.755 145.625 48.795 145.795 ;
        RECT 47.755 145.035 48.795 145.205 ;
        RECT 47.370 144.415 47.540 144.915 ;
        RECT 49.010 144.415 49.180 144.915 ;
        RECT 47.755 144.125 48.795 144.295 ;
        RECT 47.755 143.535 48.795 143.705 ;
        RECT 47.370 142.915 47.540 143.415 ;
        RECT 49.010 142.915 49.180 143.415 ;
        RECT 47.755 142.625 48.795 142.795 ;
        RECT 47.755 142.035 48.795 142.205 ;
        RECT 47.370 141.415 47.540 141.915 ;
        RECT 49.010 141.415 49.180 141.915 ;
        RECT 47.755 141.125 48.795 141.295 ;
        RECT 47.755 140.535 48.795 140.705 ;
        RECT 47.370 139.915 47.540 140.415 ;
        RECT 49.010 139.915 49.180 140.415 ;
        RECT 47.755 139.625 48.795 139.795 ;
        RECT 47.755 139.035 48.795 139.205 ;
        RECT 47.370 138.415 47.540 138.915 ;
        RECT 49.010 138.415 49.180 138.915 ;
        RECT 47.755 138.125 48.795 138.295 ;
        RECT 47.755 137.535 48.795 137.705 ;
        RECT 47.370 136.915 47.540 137.415 ;
        RECT 49.010 136.915 49.180 137.415 ;
        RECT 47.755 136.625 48.795 136.795 ;
        RECT 47.755 136.035 48.795 136.205 ;
        RECT 47.370 135.415 47.540 135.915 ;
        RECT 49.010 135.415 49.180 135.915 ;
        RECT 47.755 135.125 48.795 135.295 ;
        RECT 47.755 134.535 48.795 134.705 ;
        RECT 47.370 133.915 47.540 134.415 ;
        RECT 49.010 133.915 49.180 134.415 ;
        RECT 47.755 133.625 48.795 133.795 ;
        RECT 49.430 133.235 49.600 147.095 ;
        RECT 46.950 133.065 49.600 133.235 ;
        RECT 50.480 147.245 52.780 147.415 ;
        RECT 50.480 133.135 50.650 147.245 ;
        RECT 51.285 146.535 51.975 146.705 ;
        RECT 50.945 145.915 51.115 146.415 ;
        RECT 52.145 145.915 52.315 146.415 ;
        RECT 51.285 145.625 51.975 145.795 ;
        RECT 51.285 145.035 51.975 145.205 ;
        RECT 50.945 144.415 51.115 144.915 ;
        RECT 52.145 144.415 52.315 144.915 ;
        RECT 51.285 144.125 51.975 144.295 ;
        RECT 51.285 143.535 51.975 143.705 ;
        RECT 50.945 142.915 51.115 143.415 ;
        RECT 52.145 142.915 52.315 143.415 ;
        RECT 51.285 142.625 51.975 142.795 ;
        RECT 51.285 142.035 51.975 142.205 ;
        RECT 50.945 141.415 51.115 141.915 ;
        RECT 52.145 141.415 52.315 141.915 ;
        RECT 51.285 141.125 51.975 141.295 ;
        RECT 51.285 140.535 51.975 140.705 ;
        RECT 50.945 139.915 51.115 140.415 ;
        RECT 52.145 139.915 52.315 140.415 ;
        RECT 51.285 139.625 51.975 139.795 ;
        RECT 51.285 139.035 51.975 139.205 ;
        RECT 50.945 138.415 51.115 138.915 ;
        RECT 52.145 138.415 52.315 138.915 ;
        RECT 51.285 138.125 51.975 138.295 ;
        RECT 51.285 137.535 51.975 137.705 ;
        RECT 50.945 136.915 51.115 137.415 ;
        RECT 52.145 136.915 52.315 137.415 ;
        RECT 51.285 136.625 51.975 136.795 ;
        RECT 51.285 136.035 51.975 136.205 ;
        RECT 50.945 135.415 51.115 135.915 ;
        RECT 52.145 135.415 52.315 135.915 ;
        RECT 51.285 135.125 51.975 135.295 ;
        RECT 51.285 134.535 51.975 134.705 ;
        RECT 50.945 133.915 51.115 134.415 ;
        RECT 52.145 133.915 52.315 134.415 ;
        RECT 51.285 133.625 51.975 133.795 ;
        RECT 52.610 133.135 52.780 147.245 ;
        RECT 50.480 132.965 52.780 133.135 ;
        RECT 53.660 147.095 56.310 147.265 ;
        RECT 53.660 133.235 53.830 147.095 ;
        RECT 54.465 146.535 55.505 146.705 ;
        RECT 54.080 145.915 54.250 146.415 ;
        RECT 55.720 145.915 55.890 146.415 ;
        RECT 54.465 145.625 55.505 145.795 ;
        RECT 54.465 145.035 55.505 145.205 ;
        RECT 54.080 144.415 54.250 144.915 ;
        RECT 55.720 144.415 55.890 144.915 ;
        RECT 54.465 144.125 55.505 144.295 ;
        RECT 54.465 143.535 55.505 143.705 ;
        RECT 54.080 142.915 54.250 143.415 ;
        RECT 55.720 142.915 55.890 143.415 ;
        RECT 54.465 142.625 55.505 142.795 ;
        RECT 54.465 142.035 55.505 142.205 ;
        RECT 54.080 141.415 54.250 141.915 ;
        RECT 55.720 141.415 55.890 141.915 ;
        RECT 54.465 141.125 55.505 141.295 ;
        RECT 54.465 140.535 55.505 140.705 ;
        RECT 54.080 139.915 54.250 140.415 ;
        RECT 55.720 139.915 55.890 140.415 ;
        RECT 54.465 139.625 55.505 139.795 ;
        RECT 54.465 139.035 55.505 139.205 ;
        RECT 54.080 138.415 54.250 138.915 ;
        RECT 55.720 138.415 55.890 138.915 ;
        RECT 54.465 138.125 55.505 138.295 ;
        RECT 54.465 137.535 55.505 137.705 ;
        RECT 54.080 136.915 54.250 137.415 ;
        RECT 55.720 136.915 55.890 137.415 ;
        RECT 54.465 136.625 55.505 136.795 ;
        RECT 54.465 136.035 55.505 136.205 ;
        RECT 54.080 135.415 54.250 135.915 ;
        RECT 55.720 135.415 55.890 135.915 ;
        RECT 54.465 135.125 55.505 135.295 ;
        RECT 54.465 134.535 55.505 134.705 ;
        RECT 54.080 133.915 54.250 134.415 ;
        RECT 55.720 133.915 55.890 134.415 ;
        RECT 54.465 133.625 55.505 133.795 ;
        RECT 56.140 133.235 56.310 147.095 ;
        RECT 53.660 133.065 56.310 133.235 ;
        RECT 57.190 147.245 59.490 147.415 ;
        RECT 57.190 133.135 57.360 147.245 ;
        RECT 57.995 146.535 58.685 146.705 ;
        RECT 57.655 145.915 57.825 146.415 ;
        RECT 58.855 145.915 59.025 146.415 ;
        RECT 57.995 145.625 58.685 145.795 ;
        RECT 57.995 145.035 58.685 145.205 ;
        RECT 57.655 144.415 57.825 144.915 ;
        RECT 58.855 144.415 59.025 144.915 ;
        RECT 57.995 144.125 58.685 144.295 ;
        RECT 57.995 143.535 58.685 143.705 ;
        RECT 57.655 142.915 57.825 143.415 ;
        RECT 58.855 142.915 59.025 143.415 ;
        RECT 57.995 142.625 58.685 142.795 ;
        RECT 57.995 142.035 58.685 142.205 ;
        RECT 57.655 141.415 57.825 141.915 ;
        RECT 58.855 141.415 59.025 141.915 ;
        RECT 57.995 141.125 58.685 141.295 ;
        RECT 57.995 140.535 58.685 140.705 ;
        RECT 57.655 139.915 57.825 140.415 ;
        RECT 58.855 139.915 59.025 140.415 ;
        RECT 57.995 139.625 58.685 139.795 ;
        RECT 57.995 139.035 58.685 139.205 ;
        RECT 57.655 138.415 57.825 138.915 ;
        RECT 58.855 138.415 59.025 138.915 ;
        RECT 57.995 138.125 58.685 138.295 ;
        RECT 57.995 137.535 58.685 137.705 ;
        RECT 57.655 136.915 57.825 137.415 ;
        RECT 58.855 136.915 59.025 137.415 ;
        RECT 57.995 136.625 58.685 136.795 ;
        RECT 57.995 136.035 58.685 136.205 ;
        RECT 57.655 135.415 57.825 135.915 ;
        RECT 58.855 135.415 59.025 135.915 ;
        RECT 57.995 135.125 58.685 135.295 ;
        RECT 57.995 134.535 58.685 134.705 ;
        RECT 57.655 133.915 57.825 134.415 ;
        RECT 58.855 133.915 59.025 134.415 ;
        RECT 57.995 133.625 58.685 133.795 ;
        RECT 59.320 133.135 59.490 147.245 ;
        RECT 57.190 132.965 59.490 133.135 ;
        RECT 60.370 147.095 63.020 147.265 ;
        RECT 60.370 133.235 60.540 147.095 ;
        RECT 61.175 146.535 62.215 146.705 ;
        RECT 60.790 145.915 60.960 146.415 ;
        RECT 62.430 145.915 62.600 146.415 ;
        RECT 61.175 145.625 62.215 145.795 ;
        RECT 61.175 145.035 62.215 145.205 ;
        RECT 60.790 144.415 60.960 144.915 ;
        RECT 62.430 144.415 62.600 144.915 ;
        RECT 61.175 144.125 62.215 144.295 ;
        RECT 61.175 143.535 62.215 143.705 ;
        RECT 60.790 142.915 60.960 143.415 ;
        RECT 62.430 142.915 62.600 143.415 ;
        RECT 61.175 142.625 62.215 142.795 ;
        RECT 61.175 142.035 62.215 142.205 ;
        RECT 60.790 141.415 60.960 141.915 ;
        RECT 62.430 141.415 62.600 141.915 ;
        RECT 61.175 141.125 62.215 141.295 ;
        RECT 61.175 140.535 62.215 140.705 ;
        RECT 60.790 139.915 60.960 140.415 ;
        RECT 62.430 139.915 62.600 140.415 ;
        RECT 61.175 139.625 62.215 139.795 ;
        RECT 61.175 139.035 62.215 139.205 ;
        RECT 60.790 138.415 60.960 138.915 ;
        RECT 62.430 138.415 62.600 138.915 ;
        RECT 61.175 138.125 62.215 138.295 ;
        RECT 61.175 137.535 62.215 137.705 ;
        RECT 60.790 136.915 60.960 137.415 ;
        RECT 62.430 136.915 62.600 137.415 ;
        RECT 61.175 136.625 62.215 136.795 ;
        RECT 61.175 136.035 62.215 136.205 ;
        RECT 60.790 135.415 60.960 135.915 ;
        RECT 62.430 135.415 62.600 135.915 ;
        RECT 61.175 135.125 62.215 135.295 ;
        RECT 61.175 134.535 62.215 134.705 ;
        RECT 60.790 133.915 60.960 134.415 ;
        RECT 62.430 133.915 62.600 134.415 ;
        RECT 61.175 133.625 62.215 133.795 ;
        RECT 62.850 133.235 63.020 147.095 ;
        RECT 60.370 133.065 63.020 133.235 ;
        RECT 63.900 147.245 66.200 147.415 ;
        RECT 63.900 133.135 64.070 147.245 ;
        RECT 64.705 146.535 65.395 146.705 ;
        RECT 64.365 145.915 64.535 146.415 ;
        RECT 65.565 145.915 65.735 146.415 ;
        RECT 64.705 145.625 65.395 145.795 ;
        RECT 64.705 145.035 65.395 145.205 ;
        RECT 64.365 144.415 64.535 144.915 ;
        RECT 65.565 144.415 65.735 144.915 ;
        RECT 64.705 144.125 65.395 144.295 ;
        RECT 64.705 143.535 65.395 143.705 ;
        RECT 64.365 142.915 64.535 143.415 ;
        RECT 65.565 142.915 65.735 143.415 ;
        RECT 64.705 142.625 65.395 142.795 ;
        RECT 64.705 142.035 65.395 142.205 ;
        RECT 64.365 141.415 64.535 141.915 ;
        RECT 65.565 141.415 65.735 141.915 ;
        RECT 64.705 141.125 65.395 141.295 ;
        RECT 64.705 140.535 65.395 140.705 ;
        RECT 64.365 139.915 64.535 140.415 ;
        RECT 65.565 139.915 65.735 140.415 ;
        RECT 64.705 139.625 65.395 139.795 ;
        RECT 64.705 139.035 65.395 139.205 ;
        RECT 64.365 138.415 64.535 138.915 ;
        RECT 65.565 138.415 65.735 138.915 ;
        RECT 64.705 138.125 65.395 138.295 ;
        RECT 64.705 137.535 65.395 137.705 ;
        RECT 64.365 136.915 64.535 137.415 ;
        RECT 65.565 136.915 65.735 137.415 ;
        RECT 64.705 136.625 65.395 136.795 ;
        RECT 64.705 136.035 65.395 136.205 ;
        RECT 64.365 135.415 64.535 135.915 ;
        RECT 65.565 135.415 65.735 135.915 ;
        RECT 64.705 135.125 65.395 135.295 ;
        RECT 64.705 134.535 65.395 134.705 ;
        RECT 64.365 133.915 64.535 134.415 ;
        RECT 65.565 133.915 65.735 134.415 ;
        RECT 64.705 133.625 65.395 133.795 ;
        RECT 66.030 133.135 66.200 147.245 ;
        RECT 63.900 132.965 66.200 133.135 ;
        RECT 67.080 147.095 69.730 147.265 ;
        RECT 67.080 133.235 67.250 147.095 ;
        RECT 67.885 146.535 68.925 146.705 ;
        RECT 67.500 145.915 67.670 146.415 ;
        RECT 69.140 145.915 69.310 146.415 ;
        RECT 67.885 145.625 68.925 145.795 ;
        RECT 67.885 145.035 68.925 145.205 ;
        RECT 67.500 144.415 67.670 144.915 ;
        RECT 69.140 144.415 69.310 144.915 ;
        RECT 67.885 144.125 68.925 144.295 ;
        RECT 67.885 143.535 68.925 143.705 ;
        RECT 67.500 142.915 67.670 143.415 ;
        RECT 69.140 142.915 69.310 143.415 ;
        RECT 67.885 142.625 68.925 142.795 ;
        RECT 67.885 142.035 68.925 142.205 ;
        RECT 67.500 141.415 67.670 141.915 ;
        RECT 69.140 141.415 69.310 141.915 ;
        RECT 67.885 141.125 68.925 141.295 ;
        RECT 67.885 140.535 68.925 140.705 ;
        RECT 67.500 139.915 67.670 140.415 ;
        RECT 69.140 139.915 69.310 140.415 ;
        RECT 67.885 139.625 68.925 139.795 ;
        RECT 67.885 139.035 68.925 139.205 ;
        RECT 67.500 138.415 67.670 138.915 ;
        RECT 69.140 138.415 69.310 138.915 ;
        RECT 67.885 138.125 68.925 138.295 ;
        RECT 67.885 137.535 68.925 137.705 ;
        RECT 67.500 136.915 67.670 137.415 ;
        RECT 69.140 136.915 69.310 137.415 ;
        RECT 67.885 136.625 68.925 136.795 ;
        RECT 67.885 136.035 68.925 136.205 ;
        RECT 67.500 135.415 67.670 135.915 ;
        RECT 69.140 135.415 69.310 135.915 ;
        RECT 67.885 135.125 68.925 135.295 ;
        RECT 67.885 134.535 68.925 134.705 ;
        RECT 67.500 133.915 67.670 134.415 ;
        RECT 69.140 133.915 69.310 134.415 ;
        RECT 67.885 133.625 68.925 133.795 ;
        RECT 69.560 133.235 69.730 147.095 ;
        RECT 67.080 133.065 69.730 133.235 ;
        RECT 70.610 147.245 72.910 147.415 ;
        RECT 70.610 133.135 70.780 147.245 ;
        RECT 71.415 146.535 72.105 146.705 ;
        RECT 71.075 145.915 71.245 146.415 ;
        RECT 72.275 145.915 72.445 146.415 ;
        RECT 71.415 145.625 72.105 145.795 ;
        RECT 71.415 145.035 72.105 145.205 ;
        RECT 71.075 144.415 71.245 144.915 ;
        RECT 72.275 144.415 72.445 144.915 ;
        RECT 71.415 144.125 72.105 144.295 ;
        RECT 71.415 143.535 72.105 143.705 ;
        RECT 71.075 142.915 71.245 143.415 ;
        RECT 72.275 142.915 72.445 143.415 ;
        RECT 71.415 142.625 72.105 142.795 ;
        RECT 71.415 142.035 72.105 142.205 ;
        RECT 71.075 141.415 71.245 141.915 ;
        RECT 72.275 141.415 72.445 141.915 ;
        RECT 71.415 141.125 72.105 141.295 ;
        RECT 71.415 140.535 72.105 140.705 ;
        RECT 71.075 139.915 71.245 140.415 ;
        RECT 72.275 139.915 72.445 140.415 ;
        RECT 71.415 139.625 72.105 139.795 ;
        RECT 71.415 139.035 72.105 139.205 ;
        RECT 71.075 138.415 71.245 138.915 ;
        RECT 72.275 138.415 72.445 138.915 ;
        RECT 71.415 138.125 72.105 138.295 ;
        RECT 71.415 137.535 72.105 137.705 ;
        RECT 71.075 136.915 71.245 137.415 ;
        RECT 72.275 136.915 72.445 137.415 ;
        RECT 71.415 136.625 72.105 136.795 ;
        RECT 71.415 136.035 72.105 136.205 ;
        RECT 71.075 135.415 71.245 135.915 ;
        RECT 72.275 135.415 72.445 135.915 ;
        RECT 71.415 135.125 72.105 135.295 ;
        RECT 71.415 134.535 72.105 134.705 ;
        RECT 71.075 133.915 71.245 134.415 ;
        RECT 72.275 133.915 72.445 134.415 ;
        RECT 71.415 133.625 72.105 133.795 ;
        RECT 72.740 133.135 72.910 147.245 ;
        RECT 70.610 132.965 72.910 133.135 ;
        RECT 73.790 147.095 76.440 147.265 ;
        RECT 73.790 133.235 73.960 147.095 ;
        RECT 74.595 146.535 75.635 146.705 ;
        RECT 74.210 145.915 74.380 146.415 ;
        RECT 75.850 145.915 76.020 146.415 ;
        RECT 74.595 145.625 75.635 145.795 ;
        RECT 74.595 145.035 75.635 145.205 ;
        RECT 74.210 144.415 74.380 144.915 ;
        RECT 75.850 144.415 76.020 144.915 ;
        RECT 74.595 144.125 75.635 144.295 ;
        RECT 74.595 143.535 75.635 143.705 ;
        RECT 74.210 142.915 74.380 143.415 ;
        RECT 75.850 142.915 76.020 143.415 ;
        RECT 74.595 142.625 75.635 142.795 ;
        RECT 74.595 142.035 75.635 142.205 ;
        RECT 74.210 141.415 74.380 141.915 ;
        RECT 75.850 141.415 76.020 141.915 ;
        RECT 74.595 141.125 75.635 141.295 ;
        RECT 74.595 140.535 75.635 140.705 ;
        RECT 74.210 139.915 74.380 140.415 ;
        RECT 75.850 139.915 76.020 140.415 ;
        RECT 74.595 139.625 75.635 139.795 ;
        RECT 74.595 139.035 75.635 139.205 ;
        RECT 74.210 138.415 74.380 138.915 ;
        RECT 75.850 138.415 76.020 138.915 ;
        RECT 74.595 138.125 75.635 138.295 ;
        RECT 74.595 137.535 75.635 137.705 ;
        RECT 74.210 136.915 74.380 137.415 ;
        RECT 75.850 136.915 76.020 137.415 ;
        RECT 74.595 136.625 75.635 136.795 ;
        RECT 74.595 136.035 75.635 136.205 ;
        RECT 74.210 135.415 74.380 135.915 ;
        RECT 75.850 135.415 76.020 135.915 ;
        RECT 74.595 135.125 75.635 135.295 ;
        RECT 74.595 134.535 75.635 134.705 ;
        RECT 74.210 133.915 74.380 134.415 ;
        RECT 75.850 133.915 76.020 134.415 ;
        RECT 74.595 133.625 75.635 133.795 ;
        RECT 76.270 133.235 76.440 147.095 ;
        RECT 73.790 133.065 76.440 133.235 ;
        RECT 77.320 147.245 79.620 147.415 ;
        RECT 77.320 133.135 77.490 147.245 ;
        RECT 78.125 146.535 78.815 146.705 ;
        RECT 77.785 145.915 77.955 146.415 ;
        RECT 78.985 145.915 79.155 146.415 ;
        RECT 78.125 145.625 78.815 145.795 ;
        RECT 78.125 145.035 78.815 145.205 ;
        RECT 77.785 144.415 77.955 144.915 ;
        RECT 78.985 144.415 79.155 144.915 ;
        RECT 78.125 144.125 78.815 144.295 ;
        RECT 78.125 143.535 78.815 143.705 ;
        RECT 77.785 142.915 77.955 143.415 ;
        RECT 78.985 142.915 79.155 143.415 ;
        RECT 78.125 142.625 78.815 142.795 ;
        RECT 78.125 142.035 78.815 142.205 ;
        RECT 77.785 141.415 77.955 141.915 ;
        RECT 78.985 141.415 79.155 141.915 ;
        RECT 78.125 141.125 78.815 141.295 ;
        RECT 78.125 140.535 78.815 140.705 ;
        RECT 77.785 139.915 77.955 140.415 ;
        RECT 78.985 139.915 79.155 140.415 ;
        RECT 78.125 139.625 78.815 139.795 ;
        RECT 78.125 139.035 78.815 139.205 ;
        RECT 77.785 138.415 77.955 138.915 ;
        RECT 78.985 138.415 79.155 138.915 ;
        RECT 78.125 138.125 78.815 138.295 ;
        RECT 78.125 137.535 78.815 137.705 ;
        RECT 77.785 136.915 77.955 137.415 ;
        RECT 78.985 136.915 79.155 137.415 ;
        RECT 78.125 136.625 78.815 136.795 ;
        RECT 78.125 136.035 78.815 136.205 ;
        RECT 77.785 135.415 77.955 135.915 ;
        RECT 78.985 135.415 79.155 135.915 ;
        RECT 78.125 135.125 78.815 135.295 ;
        RECT 78.125 134.535 78.815 134.705 ;
        RECT 77.785 133.915 77.955 134.415 ;
        RECT 78.985 133.915 79.155 134.415 ;
        RECT 78.125 133.625 78.815 133.795 ;
        RECT 79.450 133.135 79.620 147.245 ;
        RECT 77.320 132.965 79.620 133.135 ;
        RECT 80.500 147.095 83.150 147.265 ;
        RECT 80.500 133.235 80.670 147.095 ;
        RECT 81.305 146.535 82.345 146.705 ;
        RECT 80.920 145.915 81.090 146.415 ;
        RECT 82.560 145.915 82.730 146.415 ;
        RECT 81.305 145.625 82.345 145.795 ;
        RECT 81.305 145.035 82.345 145.205 ;
        RECT 80.920 144.415 81.090 144.915 ;
        RECT 82.560 144.415 82.730 144.915 ;
        RECT 81.305 144.125 82.345 144.295 ;
        RECT 81.305 143.535 82.345 143.705 ;
        RECT 80.920 142.915 81.090 143.415 ;
        RECT 82.560 142.915 82.730 143.415 ;
        RECT 81.305 142.625 82.345 142.795 ;
        RECT 81.305 142.035 82.345 142.205 ;
        RECT 80.920 141.415 81.090 141.915 ;
        RECT 82.560 141.415 82.730 141.915 ;
        RECT 81.305 141.125 82.345 141.295 ;
        RECT 81.305 140.535 82.345 140.705 ;
        RECT 80.920 139.915 81.090 140.415 ;
        RECT 82.560 139.915 82.730 140.415 ;
        RECT 81.305 139.625 82.345 139.795 ;
        RECT 81.305 139.035 82.345 139.205 ;
        RECT 80.920 138.415 81.090 138.915 ;
        RECT 82.560 138.415 82.730 138.915 ;
        RECT 81.305 138.125 82.345 138.295 ;
        RECT 81.305 137.535 82.345 137.705 ;
        RECT 80.920 136.915 81.090 137.415 ;
        RECT 82.560 136.915 82.730 137.415 ;
        RECT 81.305 136.625 82.345 136.795 ;
        RECT 81.305 136.035 82.345 136.205 ;
        RECT 80.920 135.415 81.090 135.915 ;
        RECT 82.560 135.415 82.730 135.915 ;
        RECT 81.305 135.125 82.345 135.295 ;
        RECT 81.305 134.535 82.345 134.705 ;
        RECT 80.920 133.915 81.090 134.415 ;
        RECT 82.560 133.915 82.730 134.415 ;
        RECT 81.305 133.625 82.345 133.795 ;
        RECT 82.980 133.235 83.150 147.095 ;
        RECT 80.500 133.065 83.150 133.235 ;
        RECT 84.030 147.245 86.330 147.415 ;
        RECT 84.030 133.135 84.200 147.245 ;
        RECT 84.835 146.535 85.525 146.705 ;
        RECT 84.495 145.915 84.665 146.415 ;
        RECT 85.695 145.915 85.865 146.415 ;
        RECT 84.835 145.625 85.525 145.795 ;
        RECT 84.835 145.035 85.525 145.205 ;
        RECT 84.495 144.415 84.665 144.915 ;
        RECT 85.695 144.415 85.865 144.915 ;
        RECT 84.835 144.125 85.525 144.295 ;
        RECT 84.835 143.535 85.525 143.705 ;
        RECT 84.495 142.915 84.665 143.415 ;
        RECT 85.695 142.915 85.865 143.415 ;
        RECT 84.835 142.625 85.525 142.795 ;
        RECT 84.835 142.035 85.525 142.205 ;
        RECT 84.495 141.415 84.665 141.915 ;
        RECT 85.695 141.415 85.865 141.915 ;
        RECT 84.835 141.125 85.525 141.295 ;
        RECT 84.835 140.535 85.525 140.705 ;
        RECT 84.495 139.915 84.665 140.415 ;
        RECT 85.695 139.915 85.865 140.415 ;
        RECT 84.835 139.625 85.525 139.795 ;
        RECT 84.835 139.035 85.525 139.205 ;
        RECT 84.495 138.415 84.665 138.915 ;
        RECT 85.695 138.415 85.865 138.915 ;
        RECT 84.835 138.125 85.525 138.295 ;
        RECT 84.835 137.535 85.525 137.705 ;
        RECT 84.495 136.915 84.665 137.415 ;
        RECT 85.695 136.915 85.865 137.415 ;
        RECT 84.835 136.625 85.525 136.795 ;
        RECT 84.835 136.035 85.525 136.205 ;
        RECT 84.495 135.415 84.665 135.915 ;
        RECT 85.695 135.415 85.865 135.915 ;
        RECT 84.835 135.125 85.525 135.295 ;
        RECT 84.835 134.535 85.525 134.705 ;
        RECT 84.495 133.915 84.665 134.415 ;
        RECT 85.695 133.915 85.865 134.415 ;
        RECT 84.835 133.625 85.525 133.795 ;
        RECT 86.160 133.135 86.330 147.245 ;
        RECT 84.030 132.965 86.330 133.135 ;
        RECT 87.210 147.095 89.860 147.265 ;
        RECT 87.210 133.235 87.380 147.095 ;
        RECT 88.015 146.535 89.055 146.705 ;
        RECT 87.630 145.915 87.800 146.415 ;
        RECT 89.270 145.915 89.440 146.415 ;
        RECT 88.015 145.625 89.055 145.795 ;
        RECT 88.015 145.035 89.055 145.205 ;
        RECT 87.630 144.415 87.800 144.915 ;
        RECT 89.270 144.415 89.440 144.915 ;
        RECT 88.015 144.125 89.055 144.295 ;
        RECT 88.015 143.535 89.055 143.705 ;
        RECT 87.630 142.915 87.800 143.415 ;
        RECT 89.270 142.915 89.440 143.415 ;
        RECT 88.015 142.625 89.055 142.795 ;
        RECT 88.015 142.035 89.055 142.205 ;
        RECT 87.630 141.415 87.800 141.915 ;
        RECT 89.270 141.415 89.440 141.915 ;
        RECT 88.015 141.125 89.055 141.295 ;
        RECT 88.015 140.535 89.055 140.705 ;
        RECT 87.630 139.915 87.800 140.415 ;
        RECT 89.270 139.915 89.440 140.415 ;
        RECT 88.015 139.625 89.055 139.795 ;
        RECT 88.015 139.035 89.055 139.205 ;
        RECT 87.630 138.415 87.800 138.915 ;
        RECT 89.270 138.415 89.440 138.915 ;
        RECT 88.015 138.125 89.055 138.295 ;
        RECT 88.015 137.535 89.055 137.705 ;
        RECT 87.630 136.915 87.800 137.415 ;
        RECT 89.270 136.915 89.440 137.415 ;
        RECT 88.015 136.625 89.055 136.795 ;
        RECT 88.015 136.035 89.055 136.205 ;
        RECT 87.630 135.415 87.800 135.915 ;
        RECT 89.270 135.415 89.440 135.915 ;
        RECT 88.015 135.125 89.055 135.295 ;
        RECT 88.015 134.535 89.055 134.705 ;
        RECT 87.630 133.915 87.800 134.415 ;
        RECT 89.270 133.915 89.440 134.415 ;
        RECT 88.015 133.625 89.055 133.795 ;
        RECT 89.690 133.235 89.860 147.095 ;
        RECT 87.210 133.065 89.860 133.235 ;
        RECT 90.740 147.245 93.040 147.415 ;
        RECT 90.740 133.135 90.910 147.245 ;
        RECT 91.545 146.535 92.235 146.705 ;
        RECT 91.205 145.915 91.375 146.415 ;
        RECT 92.405 145.915 92.575 146.415 ;
        RECT 91.545 145.625 92.235 145.795 ;
        RECT 91.545 145.035 92.235 145.205 ;
        RECT 91.205 144.415 91.375 144.915 ;
        RECT 92.405 144.415 92.575 144.915 ;
        RECT 91.545 144.125 92.235 144.295 ;
        RECT 91.545 143.535 92.235 143.705 ;
        RECT 91.205 142.915 91.375 143.415 ;
        RECT 92.405 142.915 92.575 143.415 ;
        RECT 91.545 142.625 92.235 142.795 ;
        RECT 91.545 142.035 92.235 142.205 ;
        RECT 91.205 141.415 91.375 141.915 ;
        RECT 92.405 141.415 92.575 141.915 ;
        RECT 91.545 141.125 92.235 141.295 ;
        RECT 91.545 140.535 92.235 140.705 ;
        RECT 91.205 139.915 91.375 140.415 ;
        RECT 92.405 139.915 92.575 140.415 ;
        RECT 91.545 139.625 92.235 139.795 ;
        RECT 91.545 139.035 92.235 139.205 ;
        RECT 91.205 138.415 91.375 138.915 ;
        RECT 92.405 138.415 92.575 138.915 ;
        RECT 91.545 138.125 92.235 138.295 ;
        RECT 91.545 137.535 92.235 137.705 ;
        RECT 91.205 136.915 91.375 137.415 ;
        RECT 92.405 136.915 92.575 137.415 ;
        RECT 91.545 136.625 92.235 136.795 ;
        RECT 91.545 136.035 92.235 136.205 ;
        RECT 91.205 135.415 91.375 135.915 ;
        RECT 92.405 135.415 92.575 135.915 ;
        RECT 91.545 135.125 92.235 135.295 ;
        RECT 91.545 134.535 92.235 134.705 ;
        RECT 91.205 133.915 91.375 134.415 ;
        RECT 92.405 133.915 92.575 134.415 ;
        RECT 91.545 133.625 92.235 133.795 ;
        RECT 92.870 133.135 93.040 147.245 ;
        RECT 90.740 132.965 93.040 133.135 ;
        RECT 94.900 129.700 95.070 150.630 ;
        RECT 23.285 129.530 95.070 129.700 ;
        RECT 29.585 104.115 73.135 104.285 ;
        RECT 29.585 20.455 29.755 104.115 ;
        RECT 33.120 100.580 47.320 100.750 ;
        RECT 33.120 98.270 33.290 100.580 ;
        RECT 33.970 100.160 34.470 100.330 ;
        RECT 35.470 100.160 35.970 100.330 ;
        RECT 36.970 100.160 37.470 100.330 ;
        RECT 38.470 100.160 38.970 100.330 ;
        RECT 39.970 100.160 40.470 100.330 ;
        RECT 41.470 100.160 41.970 100.330 ;
        RECT 42.970 100.160 43.470 100.330 ;
        RECT 44.470 100.160 44.970 100.330 ;
        RECT 45.970 100.160 46.470 100.330 ;
        RECT 33.680 98.905 33.850 99.945 ;
        RECT 34.590 98.905 34.760 99.945 ;
        RECT 35.180 98.905 35.350 99.945 ;
        RECT 36.090 98.905 36.260 99.945 ;
        RECT 36.680 98.905 36.850 99.945 ;
        RECT 37.590 98.905 37.760 99.945 ;
        RECT 38.180 98.905 38.350 99.945 ;
        RECT 39.090 98.905 39.260 99.945 ;
        RECT 39.680 98.905 39.850 99.945 ;
        RECT 40.590 98.905 40.760 99.945 ;
        RECT 41.180 98.905 41.350 99.945 ;
        RECT 42.090 98.905 42.260 99.945 ;
        RECT 42.680 98.905 42.850 99.945 ;
        RECT 43.590 98.905 43.760 99.945 ;
        RECT 44.180 98.905 44.350 99.945 ;
        RECT 45.090 98.905 45.260 99.945 ;
        RECT 45.680 98.905 45.850 99.945 ;
        RECT 46.590 98.905 46.760 99.945 ;
        RECT 33.970 98.520 34.470 98.690 ;
        RECT 35.470 98.520 35.970 98.690 ;
        RECT 36.970 98.520 37.470 98.690 ;
        RECT 38.470 98.520 38.970 98.690 ;
        RECT 39.970 98.520 40.470 98.690 ;
        RECT 41.470 98.520 41.970 98.690 ;
        RECT 42.970 98.520 43.470 98.690 ;
        RECT 44.470 98.520 44.970 98.690 ;
        RECT 45.970 98.520 46.470 98.690 ;
        RECT 47.150 98.270 47.320 100.580 ;
        RECT 33.120 98.100 47.320 98.270 ;
        RECT 33.020 97.050 47.470 97.220 ;
        RECT 33.020 95.090 33.190 97.050 ;
        RECT 33.970 96.585 34.470 96.755 ;
        RECT 35.470 96.585 35.970 96.755 ;
        RECT 36.970 96.585 37.470 96.755 ;
        RECT 38.470 96.585 38.970 96.755 ;
        RECT 39.970 96.585 40.470 96.755 ;
        RECT 41.470 96.585 41.970 96.755 ;
        RECT 42.970 96.585 43.470 96.755 ;
        RECT 44.470 96.585 44.970 96.755 ;
        RECT 45.970 96.585 46.470 96.755 ;
        RECT 33.680 95.725 33.850 96.415 ;
        RECT 34.590 95.725 34.760 96.415 ;
        RECT 35.180 95.725 35.350 96.415 ;
        RECT 36.090 95.725 36.260 96.415 ;
        RECT 36.680 95.725 36.850 96.415 ;
        RECT 37.590 95.725 37.760 96.415 ;
        RECT 38.180 95.725 38.350 96.415 ;
        RECT 39.090 95.725 39.260 96.415 ;
        RECT 39.680 95.725 39.850 96.415 ;
        RECT 40.590 95.725 40.760 96.415 ;
        RECT 41.180 95.725 41.350 96.415 ;
        RECT 42.090 95.725 42.260 96.415 ;
        RECT 42.680 95.725 42.850 96.415 ;
        RECT 43.590 95.725 43.760 96.415 ;
        RECT 44.180 95.725 44.350 96.415 ;
        RECT 45.090 95.725 45.260 96.415 ;
        RECT 45.680 95.725 45.850 96.415 ;
        RECT 46.590 95.725 46.760 96.415 ;
        RECT 33.970 95.385 34.470 95.555 ;
        RECT 35.470 95.385 35.970 95.555 ;
        RECT 36.970 95.385 37.470 95.555 ;
        RECT 38.470 95.385 38.970 95.555 ;
        RECT 39.970 95.385 40.470 95.555 ;
        RECT 41.470 95.385 41.970 95.555 ;
        RECT 42.970 95.385 43.470 95.555 ;
        RECT 44.470 95.385 44.970 95.555 ;
        RECT 45.970 95.385 46.470 95.555 ;
        RECT 47.300 95.090 47.470 97.050 ;
        RECT 33.020 94.920 47.470 95.090 ;
        RECT 55.095 95.860 69.595 96.030 ;
        RECT 33.120 93.870 47.320 94.040 ;
        RECT 33.120 91.560 33.290 93.870 ;
        RECT 33.970 93.450 34.470 93.620 ;
        RECT 35.470 93.450 35.970 93.620 ;
        RECT 36.970 93.450 37.470 93.620 ;
        RECT 38.470 93.450 38.970 93.620 ;
        RECT 39.970 93.450 40.470 93.620 ;
        RECT 41.470 93.450 41.970 93.620 ;
        RECT 42.970 93.450 43.470 93.620 ;
        RECT 44.470 93.450 44.970 93.620 ;
        RECT 45.970 93.450 46.470 93.620 ;
        RECT 33.680 92.195 33.850 93.235 ;
        RECT 34.590 92.195 34.760 93.235 ;
        RECT 35.180 92.195 35.350 93.235 ;
        RECT 36.090 92.195 36.260 93.235 ;
        RECT 36.680 92.195 36.850 93.235 ;
        RECT 37.590 92.195 37.760 93.235 ;
        RECT 38.180 92.195 38.350 93.235 ;
        RECT 39.090 92.195 39.260 93.235 ;
        RECT 39.680 92.195 39.850 93.235 ;
        RECT 40.590 92.195 40.760 93.235 ;
        RECT 41.180 92.195 41.350 93.235 ;
        RECT 42.090 92.195 42.260 93.235 ;
        RECT 42.680 92.195 42.850 93.235 ;
        RECT 43.590 92.195 43.760 93.235 ;
        RECT 44.180 92.195 44.350 93.235 ;
        RECT 45.090 92.195 45.260 93.235 ;
        RECT 45.680 92.195 45.850 93.235 ;
        RECT 46.590 92.195 46.760 93.235 ;
        RECT 33.970 91.810 34.470 91.980 ;
        RECT 35.470 91.810 35.970 91.980 ;
        RECT 36.970 91.810 37.470 91.980 ;
        RECT 38.470 91.810 38.970 91.980 ;
        RECT 39.970 91.810 40.470 91.980 ;
        RECT 41.470 91.810 41.970 91.980 ;
        RECT 42.970 91.810 43.470 91.980 ;
        RECT 44.470 91.810 44.970 91.980 ;
        RECT 45.970 91.810 46.470 91.980 ;
        RECT 47.150 91.560 47.320 93.870 ;
        RECT 33.120 91.390 47.320 91.560 ;
        RECT 55.095 91.370 55.265 95.860 ;
        RECT 55.885 95.440 56.385 95.610 ;
        RECT 57.265 95.440 57.765 95.610 ;
        RECT 58.645 95.440 59.145 95.610 ;
        RECT 60.025 95.440 60.525 95.610 ;
        RECT 61.405 95.440 61.905 95.610 ;
        RECT 62.785 95.440 63.285 95.610 ;
        RECT 64.165 95.440 64.665 95.610 ;
        RECT 65.545 95.440 66.045 95.610 ;
        RECT 66.925 95.440 67.425 95.610 ;
        RECT 68.305 95.440 68.805 95.610 ;
        RECT 55.655 94.185 55.825 95.225 ;
        RECT 56.445 94.185 56.615 95.225 ;
        RECT 57.035 94.185 57.205 95.225 ;
        RECT 57.825 94.185 57.995 95.225 ;
        RECT 58.415 94.185 58.585 95.225 ;
        RECT 59.205 94.185 59.375 95.225 ;
        RECT 59.795 94.185 59.965 95.225 ;
        RECT 60.585 94.185 60.755 95.225 ;
        RECT 61.175 94.185 61.345 95.225 ;
        RECT 61.965 94.185 62.135 95.225 ;
        RECT 62.555 94.185 62.725 95.225 ;
        RECT 63.345 94.185 63.515 95.225 ;
        RECT 63.935 94.185 64.105 95.225 ;
        RECT 64.725 94.185 64.895 95.225 ;
        RECT 65.315 94.185 65.485 95.225 ;
        RECT 66.105 94.185 66.275 95.225 ;
        RECT 66.695 94.185 66.865 95.225 ;
        RECT 67.485 94.185 67.655 95.225 ;
        RECT 68.075 94.185 68.245 95.225 ;
        RECT 68.865 94.185 69.035 95.225 ;
        RECT 55.885 93.800 56.385 93.970 ;
        RECT 57.265 93.800 57.765 93.970 ;
        RECT 58.645 93.800 59.145 93.970 ;
        RECT 60.025 93.800 60.525 93.970 ;
        RECT 61.405 93.800 61.905 93.970 ;
        RECT 62.785 93.800 63.285 93.970 ;
        RECT 64.165 93.800 64.665 93.970 ;
        RECT 65.545 93.800 66.045 93.970 ;
        RECT 66.925 93.800 67.425 93.970 ;
        RECT 68.305 93.800 68.805 93.970 ;
        RECT 55.885 93.260 56.385 93.430 ;
        RECT 57.265 93.260 57.765 93.430 ;
        RECT 58.645 93.260 59.145 93.430 ;
        RECT 60.025 93.260 60.525 93.430 ;
        RECT 61.405 93.260 61.905 93.430 ;
        RECT 62.785 93.260 63.285 93.430 ;
        RECT 64.165 93.260 64.665 93.430 ;
        RECT 65.545 93.260 66.045 93.430 ;
        RECT 66.925 93.260 67.425 93.430 ;
        RECT 68.305 93.260 68.805 93.430 ;
        RECT 55.655 92.005 55.825 93.045 ;
        RECT 56.445 92.005 56.615 93.045 ;
        RECT 57.035 92.005 57.205 93.045 ;
        RECT 57.825 92.005 57.995 93.045 ;
        RECT 58.415 92.005 58.585 93.045 ;
        RECT 59.205 92.005 59.375 93.045 ;
        RECT 59.795 92.005 59.965 93.045 ;
        RECT 60.585 92.005 60.755 93.045 ;
        RECT 61.175 92.005 61.345 93.045 ;
        RECT 61.965 92.005 62.135 93.045 ;
        RECT 62.555 92.005 62.725 93.045 ;
        RECT 63.345 92.005 63.515 93.045 ;
        RECT 63.935 92.005 64.105 93.045 ;
        RECT 64.725 92.005 64.895 93.045 ;
        RECT 65.315 92.005 65.485 93.045 ;
        RECT 66.105 92.005 66.275 93.045 ;
        RECT 66.695 92.005 66.865 93.045 ;
        RECT 67.485 92.005 67.655 93.045 ;
        RECT 68.075 92.005 68.245 93.045 ;
        RECT 68.865 92.005 69.035 93.045 ;
        RECT 55.885 91.620 56.385 91.790 ;
        RECT 57.265 91.620 57.765 91.790 ;
        RECT 58.645 91.620 59.145 91.790 ;
        RECT 60.025 91.620 60.525 91.790 ;
        RECT 61.405 91.620 61.905 91.790 ;
        RECT 62.785 91.620 63.285 91.790 ;
        RECT 64.165 91.620 64.665 91.790 ;
        RECT 65.545 91.620 66.045 91.790 ;
        RECT 66.925 91.620 67.425 91.790 ;
        RECT 68.305 91.620 68.805 91.790 ;
        RECT 69.425 91.370 69.595 95.860 ;
        RECT 55.095 91.200 69.595 91.370 ;
        RECT 33.020 90.340 47.470 90.510 ;
        RECT 33.020 88.380 33.190 90.340 ;
        RECT 33.970 89.875 34.470 90.045 ;
        RECT 35.470 89.875 35.970 90.045 ;
        RECT 36.970 89.875 37.470 90.045 ;
        RECT 38.470 89.875 38.970 90.045 ;
        RECT 39.970 89.875 40.470 90.045 ;
        RECT 41.470 89.875 41.970 90.045 ;
        RECT 42.970 89.875 43.470 90.045 ;
        RECT 44.470 89.875 44.970 90.045 ;
        RECT 45.970 89.875 46.470 90.045 ;
        RECT 33.680 89.015 33.850 89.705 ;
        RECT 34.590 89.015 34.760 89.705 ;
        RECT 35.180 89.015 35.350 89.705 ;
        RECT 36.090 89.015 36.260 89.705 ;
        RECT 36.680 89.015 36.850 89.705 ;
        RECT 37.590 89.015 37.760 89.705 ;
        RECT 38.180 89.015 38.350 89.705 ;
        RECT 39.090 89.015 39.260 89.705 ;
        RECT 39.680 89.015 39.850 89.705 ;
        RECT 40.590 89.015 40.760 89.705 ;
        RECT 41.180 89.015 41.350 89.705 ;
        RECT 42.090 89.015 42.260 89.705 ;
        RECT 42.680 89.015 42.850 89.705 ;
        RECT 43.590 89.015 43.760 89.705 ;
        RECT 44.180 89.015 44.350 89.705 ;
        RECT 45.090 89.015 45.260 89.705 ;
        RECT 45.680 89.015 45.850 89.705 ;
        RECT 46.590 89.015 46.760 89.705 ;
        RECT 33.970 88.675 34.470 88.845 ;
        RECT 35.470 88.675 35.970 88.845 ;
        RECT 36.970 88.675 37.470 88.845 ;
        RECT 38.470 88.675 38.970 88.845 ;
        RECT 39.970 88.675 40.470 88.845 ;
        RECT 41.470 88.675 41.970 88.845 ;
        RECT 42.970 88.675 43.470 88.845 ;
        RECT 44.470 88.675 44.970 88.845 ;
        RECT 45.970 88.675 46.470 88.845 ;
        RECT 47.300 88.380 47.470 90.340 ;
        RECT 33.020 88.210 47.470 88.380 ;
        RECT 54.945 90.150 69.695 90.320 ;
        RECT 33.120 87.160 47.320 87.330 ;
        RECT 33.120 84.850 33.290 87.160 ;
        RECT 33.970 86.740 34.470 86.910 ;
        RECT 35.470 86.740 35.970 86.910 ;
        RECT 36.970 86.740 37.470 86.910 ;
        RECT 38.470 86.740 38.970 86.910 ;
        RECT 39.970 86.740 40.470 86.910 ;
        RECT 41.470 86.740 41.970 86.910 ;
        RECT 42.970 86.740 43.470 86.910 ;
        RECT 44.470 86.740 44.970 86.910 ;
        RECT 45.970 86.740 46.470 86.910 ;
        RECT 33.680 85.485 33.850 86.525 ;
        RECT 34.590 85.485 34.760 86.525 ;
        RECT 35.180 85.485 35.350 86.525 ;
        RECT 36.090 85.485 36.260 86.525 ;
        RECT 36.680 85.485 36.850 86.525 ;
        RECT 37.590 85.485 37.760 86.525 ;
        RECT 38.180 85.485 38.350 86.525 ;
        RECT 39.090 85.485 39.260 86.525 ;
        RECT 39.680 85.485 39.850 86.525 ;
        RECT 40.590 85.485 40.760 86.525 ;
        RECT 41.180 85.485 41.350 86.525 ;
        RECT 42.090 85.485 42.260 86.525 ;
        RECT 42.680 85.485 42.850 86.525 ;
        RECT 43.590 85.485 43.760 86.525 ;
        RECT 44.180 85.485 44.350 86.525 ;
        RECT 45.090 85.485 45.260 86.525 ;
        RECT 45.680 85.485 45.850 86.525 ;
        RECT 46.590 85.485 46.760 86.525 ;
        RECT 33.970 85.100 34.470 85.270 ;
        RECT 35.470 85.100 35.970 85.270 ;
        RECT 36.970 85.100 37.470 85.270 ;
        RECT 38.470 85.100 38.970 85.270 ;
        RECT 39.970 85.100 40.470 85.270 ;
        RECT 41.470 85.100 41.970 85.270 ;
        RECT 42.970 85.100 43.470 85.270 ;
        RECT 44.470 85.100 44.970 85.270 ;
        RECT 45.970 85.100 46.470 85.270 ;
        RECT 47.150 84.850 47.320 87.160 ;
        RECT 54.945 86.450 55.115 90.150 ;
        RECT 55.885 89.685 56.385 89.855 ;
        RECT 57.265 89.685 57.765 89.855 ;
        RECT 58.645 89.685 59.145 89.855 ;
        RECT 60.025 89.685 60.525 89.855 ;
        RECT 61.405 89.685 61.905 89.855 ;
        RECT 62.785 89.685 63.285 89.855 ;
        RECT 64.165 89.685 64.665 89.855 ;
        RECT 65.545 89.685 66.045 89.855 ;
        RECT 66.925 89.685 67.425 89.855 ;
        RECT 68.305 89.685 68.805 89.855 ;
        RECT 55.655 88.825 55.825 89.515 ;
        RECT 56.445 88.825 56.615 89.515 ;
        RECT 57.035 88.825 57.205 89.515 ;
        RECT 57.825 88.825 57.995 89.515 ;
        RECT 58.415 88.825 58.585 89.515 ;
        RECT 59.205 88.825 59.375 89.515 ;
        RECT 59.795 88.825 59.965 89.515 ;
        RECT 60.585 88.825 60.755 89.515 ;
        RECT 61.175 88.825 61.345 89.515 ;
        RECT 61.965 88.825 62.135 89.515 ;
        RECT 62.555 88.825 62.725 89.515 ;
        RECT 63.345 88.825 63.515 89.515 ;
        RECT 63.935 88.825 64.105 89.515 ;
        RECT 64.725 88.825 64.895 89.515 ;
        RECT 65.315 88.825 65.485 89.515 ;
        RECT 66.105 88.825 66.275 89.515 ;
        RECT 66.695 88.825 66.865 89.515 ;
        RECT 67.485 88.825 67.655 89.515 ;
        RECT 68.075 88.825 68.245 89.515 ;
        RECT 68.865 88.825 69.035 89.515 ;
        RECT 55.885 88.485 56.385 88.655 ;
        RECT 57.265 88.485 57.765 88.655 ;
        RECT 58.645 88.485 59.145 88.655 ;
        RECT 60.025 88.485 60.525 88.655 ;
        RECT 61.405 88.485 61.905 88.655 ;
        RECT 62.785 88.485 63.285 88.655 ;
        RECT 64.165 88.485 64.665 88.655 ;
        RECT 65.545 88.485 66.045 88.655 ;
        RECT 66.925 88.485 67.425 88.655 ;
        RECT 68.305 88.485 68.805 88.655 ;
        RECT 55.885 87.945 56.385 88.115 ;
        RECT 57.265 87.945 57.765 88.115 ;
        RECT 58.645 87.945 59.145 88.115 ;
        RECT 60.025 87.945 60.525 88.115 ;
        RECT 61.405 87.945 61.905 88.115 ;
        RECT 62.785 87.945 63.285 88.115 ;
        RECT 64.165 87.945 64.665 88.115 ;
        RECT 65.545 87.945 66.045 88.115 ;
        RECT 66.925 87.945 67.425 88.115 ;
        RECT 68.305 87.945 68.805 88.115 ;
        RECT 55.655 87.085 55.825 87.775 ;
        RECT 56.445 87.085 56.615 87.775 ;
        RECT 57.035 87.085 57.205 87.775 ;
        RECT 57.825 87.085 57.995 87.775 ;
        RECT 58.415 87.085 58.585 87.775 ;
        RECT 59.205 87.085 59.375 87.775 ;
        RECT 59.795 87.085 59.965 87.775 ;
        RECT 60.585 87.085 60.755 87.775 ;
        RECT 61.175 87.085 61.345 87.775 ;
        RECT 61.965 87.085 62.135 87.775 ;
        RECT 62.555 87.085 62.725 87.775 ;
        RECT 63.345 87.085 63.515 87.775 ;
        RECT 63.935 87.085 64.105 87.775 ;
        RECT 64.725 87.085 64.895 87.775 ;
        RECT 65.315 87.085 65.485 87.775 ;
        RECT 66.105 87.085 66.275 87.775 ;
        RECT 66.695 87.085 66.865 87.775 ;
        RECT 67.485 87.085 67.655 87.775 ;
        RECT 68.075 87.085 68.245 87.775 ;
        RECT 68.865 87.085 69.035 87.775 ;
        RECT 55.885 86.745 56.385 86.915 ;
        RECT 57.265 86.745 57.765 86.915 ;
        RECT 58.645 86.745 59.145 86.915 ;
        RECT 60.025 86.745 60.525 86.915 ;
        RECT 61.405 86.745 61.905 86.915 ;
        RECT 62.785 86.745 63.285 86.915 ;
        RECT 64.165 86.745 64.665 86.915 ;
        RECT 65.545 86.745 66.045 86.915 ;
        RECT 66.925 86.745 67.425 86.915 ;
        RECT 68.305 86.745 68.805 86.915 ;
        RECT 69.525 86.450 69.695 90.150 ;
        RECT 54.945 86.280 69.695 86.450 ;
        RECT 33.120 84.680 47.320 84.850 ;
        RECT 33.020 83.630 47.470 83.800 ;
        RECT 33.020 81.670 33.190 83.630 ;
        RECT 33.970 83.165 34.470 83.335 ;
        RECT 35.470 83.165 35.970 83.335 ;
        RECT 36.970 83.165 37.470 83.335 ;
        RECT 38.470 83.165 38.970 83.335 ;
        RECT 39.970 83.165 40.470 83.335 ;
        RECT 41.470 83.165 41.970 83.335 ;
        RECT 42.970 83.165 43.470 83.335 ;
        RECT 44.470 83.165 44.970 83.335 ;
        RECT 45.970 83.165 46.470 83.335 ;
        RECT 33.680 82.305 33.850 82.995 ;
        RECT 34.590 82.305 34.760 82.995 ;
        RECT 35.180 82.305 35.350 82.995 ;
        RECT 36.090 82.305 36.260 82.995 ;
        RECT 36.680 82.305 36.850 82.995 ;
        RECT 37.590 82.305 37.760 82.995 ;
        RECT 38.180 82.305 38.350 82.995 ;
        RECT 39.090 82.305 39.260 82.995 ;
        RECT 39.680 82.305 39.850 82.995 ;
        RECT 40.590 82.305 40.760 82.995 ;
        RECT 41.180 82.305 41.350 82.995 ;
        RECT 42.090 82.305 42.260 82.995 ;
        RECT 42.680 82.305 42.850 82.995 ;
        RECT 43.590 82.305 43.760 82.995 ;
        RECT 44.180 82.305 44.350 82.995 ;
        RECT 45.090 82.305 45.260 82.995 ;
        RECT 45.680 82.305 45.850 82.995 ;
        RECT 46.590 82.305 46.760 82.995 ;
        RECT 33.970 81.965 34.470 82.135 ;
        RECT 35.470 81.965 35.970 82.135 ;
        RECT 36.970 81.965 37.470 82.135 ;
        RECT 38.470 81.965 38.970 82.135 ;
        RECT 39.970 81.965 40.470 82.135 ;
        RECT 41.470 81.965 41.970 82.135 ;
        RECT 42.970 81.965 43.470 82.135 ;
        RECT 44.470 81.965 44.970 82.135 ;
        RECT 45.970 81.965 46.470 82.135 ;
        RECT 47.300 81.670 47.470 83.630 ;
        RECT 48.890 83.580 49.240 85.740 ;
        RECT 49.720 83.580 50.070 85.740 ;
        RECT 50.550 83.580 50.900 85.740 ;
        RECT 51.380 83.580 51.730 85.740 ;
        RECT 52.210 83.580 52.560 85.740 ;
        RECT 53.040 83.580 53.390 85.740 ;
        RECT 53.870 83.580 54.220 85.740 ;
        RECT 54.700 83.580 55.050 85.740 ;
        RECT 55.530 83.580 55.880 85.740 ;
        RECT 56.360 83.580 56.710 85.740 ;
        RECT 57.190 83.580 57.540 85.740 ;
        RECT 58.020 83.580 58.370 85.740 ;
        RECT 58.850 83.580 59.200 85.740 ;
        RECT 59.680 83.580 60.030 85.740 ;
        RECT 60.510 83.580 60.860 85.740 ;
        RECT 61.340 83.580 61.690 85.740 ;
        RECT 62.170 83.580 62.520 85.740 ;
        RECT 63.000 83.580 63.350 85.740 ;
        RECT 63.830 83.580 64.180 85.740 ;
        RECT 64.660 83.580 65.010 85.740 ;
        RECT 65.490 83.580 65.840 85.740 ;
        RECT 66.320 83.580 66.670 85.740 ;
        RECT 67.150 83.580 67.500 85.740 ;
        RECT 67.980 83.580 68.330 85.740 ;
        RECT 68.810 83.580 69.160 85.740 ;
        RECT 69.640 83.580 69.990 85.740 ;
        RECT 33.020 81.500 47.470 81.670 ;
        RECT 33.120 80.450 47.320 80.620 ;
        RECT 33.120 78.140 33.290 80.450 ;
        RECT 33.970 80.030 34.470 80.200 ;
        RECT 35.470 80.030 35.970 80.200 ;
        RECT 36.970 80.030 37.470 80.200 ;
        RECT 38.470 80.030 38.970 80.200 ;
        RECT 39.970 80.030 40.470 80.200 ;
        RECT 41.470 80.030 41.970 80.200 ;
        RECT 42.970 80.030 43.470 80.200 ;
        RECT 44.470 80.030 44.970 80.200 ;
        RECT 45.970 80.030 46.470 80.200 ;
        RECT 33.680 78.775 33.850 79.815 ;
        RECT 34.590 78.775 34.760 79.815 ;
        RECT 35.180 78.775 35.350 79.815 ;
        RECT 36.090 78.775 36.260 79.815 ;
        RECT 36.680 78.775 36.850 79.815 ;
        RECT 37.590 78.775 37.760 79.815 ;
        RECT 38.180 78.775 38.350 79.815 ;
        RECT 39.090 78.775 39.260 79.815 ;
        RECT 39.680 78.775 39.850 79.815 ;
        RECT 40.590 78.775 40.760 79.815 ;
        RECT 41.180 78.775 41.350 79.815 ;
        RECT 42.090 78.775 42.260 79.815 ;
        RECT 42.680 78.775 42.850 79.815 ;
        RECT 43.590 78.775 43.760 79.815 ;
        RECT 44.180 78.775 44.350 79.815 ;
        RECT 45.090 78.775 45.260 79.815 ;
        RECT 45.680 78.775 45.850 79.815 ;
        RECT 46.590 78.775 46.760 79.815 ;
        RECT 33.970 78.390 34.470 78.560 ;
        RECT 35.470 78.390 35.970 78.560 ;
        RECT 36.970 78.390 37.470 78.560 ;
        RECT 38.470 78.390 38.970 78.560 ;
        RECT 39.970 78.390 40.470 78.560 ;
        RECT 41.470 78.390 41.970 78.560 ;
        RECT 42.970 78.390 43.470 78.560 ;
        RECT 44.470 78.390 44.970 78.560 ;
        RECT 45.970 78.390 46.470 78.560 ;
        RECT 47.150 78.140 47.320 80.450 ;
        RECT 33.120 77.970 47.320 78.140 ;
        RECT 33.020 76.920 47.470 77.090 ;
        RECT 33.020 74.960 33.190 76.920 ;
        RECT 33.970 76.455 34.470 76.625 ;
        RECT 35.470 76.455 35.970 76.625 ;
        RECT 36.970 76.455 37.470 76.625 ;
        RECT 38.470 76.455 38.970 76.625 ;
        RECT 39.970 76.455 40.470 76.625 ;
        RECT 41.470 76.455 41.970 76.625 ;
        RECT 42.970 76.455 43.470 76.625 ;
        RECT 44.470 76.455 44.970 76.625 ;
        RECT 45.970 76.455 46.470 76.625 ;
        RECT 33.680 75.595 33.850 76.285 ;
        RECT 34.590 75.595 34.760 76.285 ;
        RECT 35.180 75.595 35.350 76.285 ;
        RECT 36.090 75.595 36.260 76.285 ;
        RECT 36.680 75.595 36.850 76.285 ;
        RECT 37.590 75.595 37.760 76.285 ;
        RECT 38.180 75.595 38.350 76.285 ;
        RECT 39.090 75.595 39.260 76.285 ;
        RECT 39.680 75.595 39.850 76.285 ;
        RECT 40.590 75.595 40.760 76.285 ;
        RECT 41.180 75.595 41.350 76.285 ;
        RECT 42.090 75.595 42.260 76.285 ;
        RECT 42.680 75.595 42.850 76.285 ;
        RECT 43.590 75.595 43.760 76.285 ;
        RECT 44.180 75.595 44.350 76.285 ;
        RECT 45.090 75.595 45.260 76.285 ;
        RECT 45.680 75.595 45.850 76.285 ;
        RECT 46.590 75.595 46.760 76.285 ;
        RECT 33.970 75.255 34.470 75.425 ;
        RECT 35.470 75.255 35.970 75.425 ;
        RECT 36.970 75.255 37.470 75.425 ;
        RECT 38.470 75.255 38.970 75.425 ;
        RECT 39.970 75.255 40.470 75.425 ;
        RECT 41.470 75.255 41.970 75.425 ;
        RECT 42.970 75.255 43.470 75.425 ;
        RECT 44.470 75.255 44.970 75.425 ;
        RECT 45.970 75.255 46.470 75.425 ;
        RECT 47.300 74.960 47.470 76.920 ;
        RECT 33.020 74.790 47.470 74.960 ;
        RECT 33.120 73.740 47.320 73.910 ;
        RECT 33.120 71.430 33.290 73.740 ;
        RECT 33.970 73.320 34.470 73.490 ;
        RECT 35.470 73.320 35.970 73.490 ;
        RECT 36.970 73.320 37.470 73.490 ;
        RECT 38.470 73.320 38.970 73.490 ;
        RECT 39.970 73.320 40.470 73.490 ;
        RECT 41.470 73.320 41.970 73.490 ;
        RECT 42.970 73.320 43.470 73.490 ;
        RECT 44.470 73.320 44.970 73.490 ;
        RECT 45.970 73.320 46.470 73.490 ;
        RECT 33.680 72.065 33.850 73.105 ;
        RECT 34.590 72.065 34.760 73.105 ;
        RECT 35.180 72.065 35.350 73.105 ;
        RECT 36.090 72.065 36.260 73.105 ;
        RECT 36.680 72.065 36.850 73.105 ;
        RECT 37.590 72.065 37.760 73.105 ;
        RECT 38.180 72.065 38.350 73.105 ;
        RECT 39.090 72.065 39.260 73.105 ;
        RECT 39.680 72.065 39.850 73.105 ;
        RECT 40.590 72.065 40.760 73.105 ;
        RECT 41.180 72.065 41.350 73.105 ;
        RECT 42.090 72.065 42.260 73.105 ;
        RECT 42.680 72.065 42.850 73.105 ;
        RECT 43.590 72.065 43.760 73.105 ;
        RECT 44.180 72.065 44.350 73.105 ;
        RECT 45.090 72.065 45.260 73.105 ;
        RECT 45.680 72.065 45.850 73.105 ;
        RECT 46.590 72.065 46.760 73.105 ;
        RECT 33.970 71.680 34.470 71.850 ;
        RECT 35.470 71.680 35.970 71.850 ;
        RECT 36.970 71.680 37.470 71.850 ;
        RECT 38.470 71.680 38.970 71.850 ;
        RECT 39.970 71.680 40.470 71.850 ;
        RECT 41.470 71.680 41.970 71.850 ;
        RECT 42.970 71.680 43.470 71.850 ;
        RECT 44.470 71.680 44.970 71.850 ;
        RECT 45.970 71.680 46.470 71.850 ;
        RECT 47.150 71.430 47.320 73.740 ;
        RECT 33.120 71.260 47.320 71.430 ;
        RECT 33.020 70.210 47.470 70.380 ;
        RECT 33.020 68.250 33.190 70.210 ;
        RECT 33.970 69.745 34.470 69.915 ;
        RECT 35.470 69.745 35.970 69.915 ;
        RECT 36.970 69.745 37.470 69.915 ;
        RECT 38.470 69.745 38.970 69.915 ;
        RECT 39.970 69.745 40.470 69.915 ;
        RECT 41.470 69.745 41.970 69.915 ;
        RECT 42.970 69.745 43.470 69.915 ;
        RECT 44.470 69.745 44.970 69.915 ;
        RECT 45.970 69.745 46.470 69.915 ;
        RECT 33.680 68.885 33.850 69.575 ;
        RECT 34.590 68.885 34.760 69.575 ;
        RECT 35.180 68.885 35.350 69.575 ;
        RECT 36.090 68.885 36.260 69.575 ;
        RECT 36.680 68.885 36.850 69.575 ;
        RECT 37.590 68.885 37.760 69.575 ;
        RECT 38.180 68.885 38.350 69.575 ;
        RECT 39.090 68.885 39.260 69.575 ;
        RECT 39.680 68.885 39.850 69.575 ;
        RECT 40.590 68.885 40.760 69.575 ;
        RECT 41.180 68.885 41.350 69.575 ;
        RECT 42.090 68.885 42.260 69.575 ;
        RECT 42.680 68.885 42.850 69.575 ;
        RECT 43.590 68.885 43.760 69.575 ;
        RECT 44.180 68.885 44.350 69.575 ;
        RECT 45.090 68.885 45.260 69.575 ;
        RECT 45.680 68.885 45.850 69.575 ;
        RECT 46.590 68.885 46.760 69.575 ;
        RECT 33.970 68.545 34.470 68.715 ;
        RECT 35.470 68.545 35.970 68.715 ;
        RECT 36.970 68.545 37.470 68.715 ;
        RECT 38.470 68.545 38.970 68.715 ;
        RECT 39.970 68.545 40.470 68.715 ;
        RECT 41.470 68.545 41.970 68.715 ;
        RECT 42.970 68.545 43.470 68.715 ;
        RECT 44.470 68.545 44.970 68.715 ;
        RECT 45.970 68.545 46.470 68.715 ;
        RECT 47.300 68.250 47.470 70.210 ;
        RECT 33.020 68.080 47.470 68.250 ;
        RECT 33.120 67.030 47.320 67.200 ;
        RECT 33.120 64.720 33.290 67.030 ;
        RECT 33.970 66.610 34.470 66.780 ;
        RECT 35.470 66.610 35.970 66.780 ;
        RECT 36.970 66.610 37.470 66.780 ;
        RECT 38.470 66.610 38.970 66.780 ;
        RECT 39.970 66.610 40.470 66.780 ;
        RECT 41.470 66.610 41.970 66.780 ;
        RECT 42.970 66.610 43.470 66.780 ;
        RECT 44.470 66.610 44.970 66.780 ;
        RECT 45.970 66.610 46.470 66.780 ;
        RECT 33.680 65.355 33.850 66.395 ;
        RECT 34.590 65.355 34.760 66.395 ;
        RECT 35.180 65.355 35.350 66.395 ;
        RECT 36.090 65.355 36.260 66.395 ;
        RECT 36.680 65.355 36.850 66.395 ;
        RECT 37.590 65.355 37.760 66.395 ;
        RECT 38.180 65.355 38.350 66.395 ;
        RECT 39.090 65.355 39.260 66.395 ;
        RECT 39.680 65.355 39.850 66.395 ;
        RECT 40.590 65.355 40.760 66.395 ;
        RECT 41.180 65.355 41.350 66.395 ;
        RECT 42.090 65.355 42.260 66.395 ;
        RECT 42.680 65.355 42.850 66.395 ;
        RECT 43.590 65.355 43.760 66.395 ;
        RECT 44.180 65.355 44.350 66.395 ;
        RECT 45.090 65.355 45.260 66.395 ;
        RECT 45.680 65.355 45.850 66.395 ;
        RECT 46.590 65.355 46.760 66.395 ;
        RECT 33.970 64.970 34.470 65.140 ;
        RECT 35.470 64.970 35.970 65.140 ;
        RECT 36.970 64.970 37.470 65.140 ;
        RECT 38.470 64.970 38.970 65.140 ;
        RECT 39.970 64.970 40.470 65.140 ;
        RECT 41.470 64.970 41.970 65.140 ;
        RECT 42.970 64.970 43.470 65.140 ;
        RECT 44.470 64.970 44.970 65.140 ;
        RECT 45.970 64.970 46.470 65.140 ;
        RECT 47.150 64.720 47.320 67.030 ;
        RECT 33.120 64.550 47.320 64.720 ;
        RECT 33.020 63.500 47.470 63.670 ;
        RECT 33.020 61.540 33.190 63.500 ;
        RECT 33.970 63.035 34.470 63.205 ;
        RECT 35.470 63.035 35.970 63.205 ;
        RECT 36.970 63.035 37.470 63.205 ;
        RECT 38.470 63.035 38.970 63.205 ;
        RECT 39.970 63.035 40.470 63.205 ;
        RECT 41.470 63.035 41.970 63.205 ;
        RECT 42.970 63.035 43.470 63.205 ;
        RECT 44.470 63.035 44.970 63.205 ;
        RECT 45.970 63.035 46.470 63.205 ;
        RECT 33.680 62.175 33.850 62.865 ;
        RECT 34.590 62.175 34.760 62.865 ;
        RECT 35.180 62.175 35.350 62.865 ;
        RECT 36.090 62.175 36.260 62.865 ;
        RECT 36.680 62.175 36.850 62.865 ;
        RECT 37.590 62.175 37.760 62.865 ;
        RECT 38.180 62.175 38.350 62.865 ;
        RECT 39.090 62.175 39.260 62.865 ;
        RECT 39.680 62.175 39.850 62.865 ;
        RECT 40.590 62.175 40.760 62.865 ;
        RECT 41.180 62.175 41.350 62.865 ;
        RECT 42.090 62.175 42.260 62.865 ;
        RECT 42.680 62.175 42.850 62.865 ;
        RECT 43.590 62.175 43.760 62.865 ;
        RECT 44.180 62.175 44.350 62.865 ;
        RECT 45.090 62.175 45.260 62.865 ;
        RECT 45.680 62.175 45.850 62.865 ;
        RECT 46.590 62.175 46.760 62.865 ;
        RECT 33.970 61.835 34.470 62.005 ;
        RECT 35.470 61.835 35.970 62.005 ;
        RECT 36.970 61.835 37.470 62.005 ;
        RECT 38.470 61.835 38.970 62.005 ;
        RECT 39.970 61.835 40.470 62.005 ;
        RECT 41.470 61.835 41.970 62.005 ;
        RECT 42.970 61.835 43.470 62.005 ;
        RECT 44.470 61.835 44.970 62.005 ;
        RECT 45.970 61.835 46.470 62.005 ;
        RECT 47.300 61.540 47.470 63.500 ;
        RECT 33.020 61.370 47.470 61.540 ;
        RECT 33.120 60.320 47.320 60.490 ;
        RECT 33.120 58.010 33.290 60.320 ;
        RECT 33.970 59.900 34.470 60.070 ;
        RECT 35.470 59.900 35.970 60.070 ;
        RECT 36.970 59.900 37.470 60.070 ;
        RECT 38.470 59.900 38.970 60.070 ;
        RECT 39.970 59.900 40.470 60.070 ;
        RECT 41.470 59.900 41.970 60.070 ;
        RECT 42.970 59.900 43.470 60.070 ;
        RECT 44.470 59.900 44.970 60.070 ;
        RECT 45.970 59.900 46.470 60.070 ;
        RECT 33.680 58.645 33.850 59.685 ;
        RECT 34.590 58.645 34.760 59.685 ;
        RECT 35.180 58.645 35.350 59.685 ;
        RECT 36.090 58.645 36.260 59.685 ;
        RECT 36.680 58.645 36.850 59.685 ;
        RECT 37.590 58.645 37.760 59.685 ;
        RECT 38.180 58.645 38.350 59.685 ;
        RECT 39.090 58.645 39.260 59.685 ;
        RECT 39.680 58.645 39.850 59.685 ;
        RECT 40.590 58.645 40.760 59.685 ;
        RECT 41.180 58.645 41.350 59.685 ;
        RECT 42.090 58.645 42.260 59.685 ;
        RECT 42.680 58.645 42.850 59.685 ;
        RECT 43.590 58.645 43.760 59.685 ;
        RECT 44.180 58.645 44.350 59.685 ;
        RECT 45.090 58.645 45.260 59.685 ;
        RECT 45.680 58.645 45.850 59.685 ;
        RECT 46.590 58.645 46.760 59.685 ;
        RECT 33.970 58.260 34.470 58.430 ;
        RECT 35.470 58.260 35.970 58.430 ;
        RECT 36.970 58.260 37.470 58.430 ;
        RECT 38.470 58.260 38.970 58.430 ;
        RECT 39.970 58.260 40.470 58.430 ;
        RECT 41.470 58.260 41.970 58.430 ;
        RECT 42.970 58.260 43.470 58.430 ;
        RECT 44.470 58.260 44.970 58.430 ;
        RECT 45.970 58.260 46.470 58.430 ;
        RECT 47.150 58.010 47.320 60.320 ;
        RECT 33.120 57.840 47.320 58.010 ;
        RECT 33.020 56.790 47.470 56.960 ;
        RECT 33.020 54.830 33.190 56.790 ;
        RECT 33.970 56.325 34.470 56.495 ;
        RECT 35.470 56.325 35.970 56.495 ;
        RECT 36.970 56.325 37.470 56.495 ;
        RECT 38.470 56.325 38.970 56.495 ;
        RECT 39.970 56.325 40.470 56.495 ;
        RECT 41.470 56.325 41.970 56.495 ;
        RECT 42.970 56.325 43.470 56.495 ;
        RECT 44.470 56.325 44.970 56.495 ;
        RECT 45.970 56.325 46.470 56.495 ;
        RECT 33.680 55.465 33.850 56.155 ;
        RECT 34.590 55.465 34.760 56.155 ;
        RECT 35.180 55.465 35.350 56.155 ;
        RECT 36.090 55.465 36.260 56.155 ;
        RECT 36.680 55.465 36.850 56.155 ;
        RECT 37.590 55.465 37.760 56.155 ;
        RECT 38.180 55.465 38.350 56.155 ;
        RECT 39.090 55.465 39.260 56.155 ;
        RECT 39.680 55.465 39.850 56.155 ;
        RECT 40.590 55.465 40.760 56.155 ;
        RECT 41.180 55.465 41.350 56.155 ;
        RECT 42.090 55.465 42.260 56.155 ;
        RECT 42.680 55.465 42.850 56.155 ;
        RECT 43.590 55.465 43.760 56.155 ;
        RECT 44.180 55.465 44.350 56.155 ;
        RECT 45.090 55.465 45.260 56.155 ;
        RECT 45.680 55.465 45.850 56.155 ;
        RECT 46.590 55.465 46.760 56.155 ;
        RECT 33.970 55.125 34.470 55.295 ;
        RECT 35.470 55.125 35.970 55.295 ;
        RECT 36.970 55.125 37.470 55.295 ;
        RECT 38.470 55.125 38.970 55.295 ;
        RECT 39.970 55.125 40.470 55.295 ;
        RECT 41.470 55.125 41.970 55.295 ;
        RECT 42.970 55.125 43.470 55.295 ;
        RECT 44.470 55.125 44.970 55.295 ;
        RECT 45.970 55.125 46.470 55.295 ;
        RECT 47.300 54.830 47.470 56.790 ;
        RECT 33.020 54.660 47.470 54.830 ;
        RECT 33.120 53.610 47.320 53.780 ;
        RECT 33.120 51.300 33.290 53.610 ;
        RECT 33.970 53.190 34.470 53.360 ;
        RECT 35.470 53.190 35.970 53.360 ;
        RECT 36.970 53.190 37.470 53.360 ;
        RECT 38.470 53.190 38.970 53.360 ;
        RECT 39.970 53.190 40.470 53.360 ;
        RECT 41.470 53.190 41.970 53.360 ;
        RECT 42.970 53.190 43.470 53.360 ;
        RECT 44.470 53.190 44.970 53.360 ;
        RECT 45.970 53.190 46.470 53.360 ;
        RECT 33.680 51.935 33.850 52.975 ;
        RECT 34.590 51.935 34.760 52.975 ;
        RECT 35.180 51.935 35.350 52.975 ;
        RECT 36.090 51.935 36.260 52.975 ;
        RECT 36.680 51.935 36.850 52.975 ;
        RECT 37.590 51.935 37.760 52.975 ;
        RECT 38.180 51.935 38.350 52.975 ;
        RECT 39.090 51.935 39.260 52.975 ;
        RECT 39.680 51.935 39.850 52.975 ;
        RECT 40.590 51.935 40.760 52.975 ;
        RECT 41.180 51.935 41.350 52.975 ;
        RECT 42.090 51.935 42.260 52.975 ;
        RECT 42.680 51.935 42.850 52.975 ;
        RECT 43.590 51.935 43.760 52.975 ;
        RECT 44.180 51.935 44.350 52.975 ;
        RECT 45.090 51.935 45.260 52.975 ;
        RECT 45.680 51.935 45.850 52.975 ;
        RECT 46.590 51.935 46.760 52.975 ;
        RECT 33.970 51.550 34.470 51.720 ;
        RECT 35.470 51.550 35.970 51.720 ;
        RECT 36.970 51.550 37.470 51.720 ;
        RECT 38.470 51.550 38.970 51.720 ;
        RECT 39.970 51.550 40.470 51.720 ;
        RECT 41.470 51.550 41.970 51.720 ;
        RECT 42.970 51.550 43.470 51.720 ;
        RECT 44.470 51.550 44.970 51.720 ;
        RECT 45.970 51.550 46.470 51.720 ;
        RECT 47.150 51.300 47.320 53.610 ;
        RECT 33.120 51.130 47.320 51.300 ;
        RECT 33.020 50.080 47.470 50.250 ;
        RECT 33.020 48.120 33.190 50.080 ;
        RECT 33.970 49.615 34.470 49.785 ;
        RECT 35.470 49.615 35.970 49.785 ;
        RECT 36.970 49.615 37.470 49.785 ;
        RECT 38.470 49.615 38.970 49.785 ;
        RECT 39.970 49.615 40.470 49.785 ;
        RECT 41.470 49.615 41.970 49.785 ;
        RECT 42.970 49.615 43.470 49.785 ;
        RECT 44.470 49.615 44.970 49.785 ;
        RECT 45.970 49.615 46.470 49.785 ;
        RECT 33.680 48.755 33.850 49.445 ;
        RECT 34.590 48.755 34.760 49.445 ;
        RECT 35.180 48.755 35.350 49.445 ;
        RECT 36.090 48.755 36.260 49.445 ;
        RECT 36.680 48.755 36.850 49.445 ;
        RECT 37.590 48.755 37.760 49.445 ;
        RECT 38.180 48.755 38.350 49.445 ;
        RECT 39.090 48.755 39.260 49.445 ;
        RECT 39.680 48.755 39.850 49.445 ;
        RECT 40.590 48.755 40.760 49.445 ;
        RECT 41.180 48.755 41.350 49.445 ;
        RECT 42.090 48.755 42.260 49.445 ;
        RECT 42.680 48.755 42.850 49.445 ;
        RECT 43.590 48.755 43.760 49.445 ;
        RECT 44.180 48.755 44.350 49.445 ;
        RECT 45.090 48.755 45.260 49.445 ;
        RECT 45.680 48.755 45.850 49.445 ;
        RECT 46.590 48.755 46.760 49.445 ;
        RECT 33.970 48.415 34.470 48.585 ;
        RECT 35.470 48.415 35.970 48.585 ;
        RECT 36.970 48.415 37.470 48.585 ;
        RECT 38.470 48.415 38.970 48.585 ;
        RECT 39.970 48.415 40.470 48.585 ;
        RECT 41.470 48.415 41.970 48.585 ;
        RECT 42.970 48.415 43.470 48.585 ;
        RECT 44.470 48.415 44.970 48.585 ;
        RECT 45.970 48.415 46.470 48.585 ;
        RECT 47.300 48.120 47.470 50.080 ;
        RECT 48.890 49.580 49.240 51.740 ;
        RECT 49.720 49.580 50.070 51.740 ;
        RECT 50.550 49.580 50.900 51.740 ;
        RECT 51.380 49.580 51.730 51.740 ;
        RECT 52.210 49.580 52.560 51.740 ;
        RECT 53.040 49.580 53.390 51.740 ;
        RECT 53.870 49.580 54.220 51.740 ;
        RECT 54.700 49.580 55.050 51.740 ;
        RECT 55.530 49.580 55.880 51.740 ;
        RECT 56.360 49.580 56.710 51.740 ;
        RECT 57.190 49.580 57.540 51.740 ;
        RECT 58.020 49.580 58.370 51.740 ;
        RECT 58.850 49.580 59.200 51.740 ;
        RECT 59.680 49.580 60.030 51.740 ;
        RECT 60.510 49.580 60.860 51.740 ;
        RECT 61.340 49.580 61.690 51.740 ;
        RECT 62.170 49.580 62.520 51.740 ;
        RECT 63.000 49.580 63.350 51.740 ;
        RECT 63.830 49.580 64.180 51.740 ;
        RECT 64.660 49.580 65.010 51.740 ;
        RECT 65.490 49.580 65.840 51.740 ;
        RECT 66.320 49.580 66.670 51.740 ;
        RECT 67.150 49.580 67.500 51.740 ;
        RECT 67.980 49.580 68.330 51.740 ;
        RECT 68.810 49.580 69.160 51.740 ;
        RECT 69.640 49.580 69.990 51.740 ;
        RECT 33.020 47.950 47.470 48.120 ;
        RECT 55.100 48.825 69.600 48.995 ;
        RECT 33.120 46.900 47.320 47.070 ;
        RECT 33.120 44.590 33.290 46.900 ;
        RECT 33.970 46.480 34.470 46.650 ;
        RECT 35.470 46.480 35.970 46.650 ;
        RECT 36.970 46.480 37.470 46.650 ;
        RECT 38.470 46.480 38.970 46.650 ;
        RECT 39.970 46.480 40.470 46.650 ;
        RECT 41.470 46.480 41.970 46.650 ;
        RECT 42.970 46.480 43.470 46.650 ;
        RECT 44.470 46.480 44.970 46.650 ;
        RECT 45.970 46.480 46.470 46.650 ;
        RECT 33.680 45.225 33.850 46.265 ;
        RECT 34.590 45.225 34.760 46.265 ;
        RECT 35.180 45.225 35.350 46.265 ;
        RECT 36.090 45.225 36.260 46.265 ;
        RECT 36.680 45.225 36.850 46.265 ;
        RECT 37.590 45.225 37.760 46.265 ;
        RECT 38.180 45.225 38.350 46.265 ;
        RECT 39.090 45.225 39.260 46.265 ;
        RECT 39.680 45.225 39.850 46.265 ;
        RECT 40.590 45.225 40.760 46.265 ;
        RECT 41.180 45.225 41.350 46.265 ;
        RECT 42.090 45.225 42.260 46.265 ;
        RECT 42.680 45.225 42.850 46.265 ;
        RECT 43.590 45.225 43.760 46.265 ;
        RECT 44.180 45.225 44.350 46.265 ;
        RECT 45.090 45.225 45.260 46.265 ;
        RECT 45.680 45.225 45.850 46.265 ;
        RECT 46.590 45.225 46.760 46.265 ;
        RECT 33.970 44.840 34.470 45.010 ;
        RECT 35.470 44.840 35.970 45.010 ;
        RECT 36.970 44.840 37.470 45.010 ;
        RECT 38.470 44.840 38.970 45.010 ;
        RECT 39.970 44.840 40.470 45.010 ;
        RECT 41.470 44.840 41.970 45.010 ;
        RECT 42.970 44.840 43.470 45.010 ;
        RECT 44.470 44.840 44.970 45.010 ;
        RECT 45.970 44.840 46.470 45.010 ;
        RECT 47.150 44.590 47.320 46.900 ;
        RECT 33.120 44.420 47.320 44.590 ;
        RECT 55.100 44.335 55.270 48.825 ;
        RECT 55.890 48.405 56.390 48.575 ;
        RECT 57.270 48.405 57.770 48.575 ;
        RECT 58.650 48.405 59.150 48.575 ;
        RECT 60.030 48.405 60.530 48.575 ;
        RECT 61.410 48.405 61.910 48.575 ;
        RECT 62.790 48.405 63.290 48.575 ;
        RECT 64.170 48.405 64.670 48.575 ;
        RECT 65.550 48.405 66.050 48.575 ;
        RECT 66.930 48.405 67.430 48.575 ;
        RECT 68.310 48.405 68.810 48.575 ;
        RECT 55.660 47.150 55.830 48.190 ;
        RECT 56.450 47.150 56.620 48.190 ;
        RECT 57.040 47.150 57.210 48.190 ;
        RECT 57.830 47.150 58.000 48.190 ;
        RECT 58.420 47.150 58.590 48.190 ;
        RECT 59.210 47.150 59.380 48.190 ;
        RECT 59.800 47.150 59.970 48.190 ;
        RECT 60.590 47.150 60.760 48.190 ;
        RECT 61.180 47.150 61.350 48.190 ;
        RECT 61.970 47.150 62.140 48.190 ;
        RECT 62.560 47.150 62.730 48.190 ;
        RECT 63.350 47.150 63.520 48.190 ;
        RECT 63.940 47.150 64.110 48.190 ;
        RECT 64.730 47.150 64.900 48.190 ;
        RECT 65.320 47.150 65.490 48.190 ;
        RECT 66.110 47.150 66.280 48.190 ;
        RECT 66.700 47.150 66.870 48.190 ;
        RECT 67.490 47.150 67.660 48.190 ;
        RECT 68.080 47.150 68.250 48.190 ;
        RECT 68.870 47.150 69.040 48.190 ;
        RECT 55.890 46.765 56.390 46.935 ;
        RECT 57.270 46.765 57.770 46.935 ;
        RECT 58.650 46.765 59.150 46.935 ;
        RECT 60.030 46.765 60.530 46.935 ;
        RECT 61.410 46.765 61.910 46.935 ;
        RECT 62.790 46.765 63.290 46.935 ;
        RECT 64.170 46.765 64.670 46.935 ;
        RECT 65.550 46.765 66.050 46.935 ;
        RECT 66.930 46.765 67.430 46.935 ;
        RECT 68.310 46.765 68.810 46.935 ;
        RECT 55.890 46.225 56.390 46.395 ;
        RECT 57.270 46.225 57.770 46.395 ;
        RECT 58.650 46.225 59.150 46.395 ;
        RECT 60.030 46.225 60.530 46.395 ;
        RECT 61.410 46.225 61.910 46.395 ;
        RECT 62.790 46.225 63.290 46.395 ;
        RECT 64.170 46.225 64.670 46.395 ;
        RECT 65.550 46.225 66.050 46.395 ;
        RECT 66.930 46.225 67.430 46.395 ;
        RECT 68.310 46.225 68.810 46.395 ;
        RECT 55.660 44.970 55.830 46.010 ;
        RECT 56.450 44.970 56.620 46.010 ;
        RECT 57.040 44.970 57.210 46.010 ;
        RECT 57.830 44.970 58.000 46.010 ;
        RECT 58.420 44.970 58.590 46.010 ;
        RECT 59.210 44.970 59.380 46.010 ;
        RECT 59.800 44.970 59.970 46.010 ;
        RECT 60.590 44.970 60.760 46.010 ;
        RECT 61.180 44.970 61.350 46.010 ;
        RECT 61.970 44.970 62.140 46.010 ;
        RECT 62.560 44.970 62.730 46.010 ;
        RECT 63.350 44.970 63.520 46.010 ;
        RECT 63.940 44.970 64.110 46.010 ;
        RECT 64.730 44.970 64.900 46.010 ;
        RECT 65.320 44.970 65.490 46.010 ;
        RECT 66.110 44.970 66.280 46.010 ;
        RECT 66.700 44.970 66.870 46.010 ;
        RECT 67.490 44.970 67.660 46.010 ;
        RECT 68.080 44.970 68.250 46.010 ;
        RECT 68.870 44.970 69.040 46.010 ;
        RECT 55.890 44.585 56.390 44.755 ;
        RECT 57.270 44.585 57.770 44.755 ;
        RECT 58.650 44.585 59.150 44.755 ;
        RECT 60.030 44.585 60.530 44.755 ;
        RECT 61.410 44.585 61.910 44.755 ;
        RECT 62.790 44.585 63.290 44.755 ;
        RECT 64.170 44.585 64.670 44.755 ;
        RECT 65.550 44.585 66.050 44.755 ;
        RECT 66.930 44.585 67.430 44.755 ;
        RECT 68.310 44.585 68.810 44.755 ;
        RECT 69.430 44.335 69.600 48.825 ;
        RECT 55.100 44.165 69.600 44.335 ;
        RECT 33.020 43.370 47.470 43.540 ;
        RECT 33.020 41.410 33.190 43.370 ;
        RECT 33.970 42.905 34.470 43.075 ;
        RECT 35.470 42.905 35.970 43.075 ;
        RECT 36.970 42.905 37.470 43.075 ;
        RECT 38.470 42.905 38.970 43.075 ;
        RECT 39.970 42.905 40.470 43.075 ;
        RECT 41.470 42.905 41.970 43.075 ;
        RECT 42.970 42.905 43.470 43.075 ;
        RECT 44.470 42.905 44.970 43.075 ;
        RECT 45.970 42.905 46.470 43.075 ;
        RECT 33.680 42.045 33.850 42.735 ;
        RECT 34.590 42.045 34.760 42.735 ;
        RECT 35.180 42.045 35.350 42.735 ;
        RECT 36.090 42.045 36.260 42.735 ;
        RECT 36.680 42.045 36.850 42.735 ;
        RECT 37.590 42.045 37.760 42.735 ;
        RECT 38.180 42.045 38.350 42.735 ;
        RECT 39.090 42.045 39.260 42.735 ;
        RECT 39.680 42.045 39.850 42.735 ;
        RECT 40.590 42.045 40.760 42.735 ;
        RECT 41.180 42.045 41.350 42.735 ;
        RECT 42.090 42.045 42.260 42.735 ;
        RECT 42.680 42.045 42.850 42.735 ;
        RECT 43.590 42.045 43.760 42.735 ;
        RECT 44.180 42.045 44.350 42.735 ;
        RECT 45.090 42.045 45.260 42.735 ;
        RECT 45.680 42.045 45.850 42.735 ;
        RECT 46.590 42.045 46.760 42.735 ;
        RECT 33.970 41.705 34.470 41.875 ;
        RECT 35.470 41.705 35.970 41.875 ;
        RECT 36.970 41.705 37.470 41.875 ;
        RECT 38.470 41.705 38.970 41.875 ;
        RECT 39.970 41.705 40.470 41.875 ;
        RECT 41.470 41.705 41.970 41.875 ;
        RECT 42.970 41.705 43.470 41.875 ;
        RECT 44.470 41.705 44.970 41.875 ;
        RECT 45.970 41.705 46.470 41.875 ;
        RECT 47.300 41.410 47.470 43.370 ;
        RECT 33.020 41.240 47.470 41.410 ;
        RECT 54.950 43.115 69.700 43.285 ;
        RECT 33.120 40.190 47.320 40.360 ;
        RECT 33.120 37.880 33.290 40.190 ;
        RECT 33.970 39.770 34.470 39.940 ;
        RECT 35.470 39.770 35.970 39.940 ;
        RECT 36.970 39.770 37.470 39.940 ;
        RECT 38.470 39.770 38.970 39.940 ;
        RECT 39.970 39.770 40.470 39.940 ;
        RECT 41.470 39.770 41.970 39.940 ;
        RECT 42.970 39.770 43.470 39.940 ;
        RECT 44.470 39.770 44.970 39.940 ;
        RECT 45.970 39.770 46.470 39.940 ;
        RECT 33.680 38.515 33.850 39.555 ;
        RECT 34.590 38.515 34.760 39.555 ;
        RECT 35.180 38.515 35.350 39.555 ;
        RECT 36.090 38.515 36.260 39.555 ;
        RECT 36.680 38.515 36.850 39.555 ;
        RECT 37.590 38.515 37.760 39.555 ;
        RECT 38.180 38.515 38.350 39.555 ;
        RECT 39.090 38.515 39.260 39.555 ;
        RECT 39.680 38.515 39.850 39.555 ;
        RECT 40.590 38.515 40.760 39.555 ;
        RECT 41.180 38.515 41.350 39.555 ;
        RECT 42.090 38.515 42.260 39.555 ;
        RECT 42.680 38.515 42.850 39.555 ;
        RECT 43.590 38.515 43.760 39.555 ;
        RECT 44.180 38.515 44.350 39.555 ;
        RECT 45.090 38.515 45.260 39.555 ;
        RECT 45.680 38.515 45.850 39.555 ;
        RECT 46.590 38.515 46.760 39.555 ;
        RECT 33.970 38.130 34.470 38.300 ;
        RECT 35.470 38.130 35.970 38.300 ;
        RECT 36.970 38.130 37.470 38.300 ;
        RECT 38.470 38.130 38.970 38.300 ;
        RECT 39.970 38.130 40.470 38.300 ;
        RECT 41.470 38.130 41.970 38.300 ;
        RECT 42.970 38.130 43.470 38.300 ;
        RECT 44.470 38.130 44.970 38.300 ;
        RECT 45.970 38.130 46.470 38.300 ;
        RECT 47.150 37.880 47.320 40.190 ;
        RECT 54.950 39.415 55.120 43.115 ;
        RECT 55.890 42.650 56.390 42.820 ;
        RECT 57.270 42.650 57.770 42.820 ;
        RECT 58.650 42.650 59.150 42.820 ;
        RECT 60.030 42.650 60.530 42.820 ;
        RECT 61.410 42.650 61.910 42.820 ;
        RECT 62.790 42.650 63.290 42.820 ;
        RECT 64.170 42.650 64.670 42.820 ;
        RECT 65.550 42.650 66.050 42.820 ;
        RECT 66.930 42.650 67.430 42.820 ;
        RECT 68.310 42.650 68.810 42.820 ;
        RECT 55.660 41.790 55.830 42.480 ;
        RECT 56.450 41.790 56.620 42.480 ;
        RECT 57.040 41.790 57.210 42.480 ;
        RECT 57.830 41.790 58.000 42.480 ;
        RECT 58.420 41.790 58.590 42.480 ;
        RECT 59.210 41.790 59.380 42.480 ;
        RECT 59.800 41.790 59.970 42.480 ;
        RECT 60.590 41.790 60.760 42.480 ;
        RECT 61.180 41.790 61.350 42.480 ;
        RECT 61.970 41.790 62.140 42.480 ;
        RECT 62.560 41.790 62.730 42.480 ;
        RECT 63.350 41.790 63.520 42.480 ;
        RECT 63.940 41.790 64.110 42.480 ;
        RECT 64.730 41.790 64.900 42.480 ;
        RECT 65.320 41.790 65.490 42.480 ;
        RECT 66.110 41.790 66.280 42.480 ;
        RECT 66.700 41.790 66.870 42.480 ;
        RECT 67.490 41.790 67.660 42.480 ;
        RECT 68.080 41.790 68.250 42.480 ;
        RECT 68.870 41.790 69.040 42.480 ;
        RECT 55.890 41.450 56.390 41.620 ;
        RECT 57.270 41.450 57.770 41.620 ;
        RECT 58.650 41.450 59.150 41.620 ;
        RECT 60.030 41.450 60.530 41.620 ;
        RECT 61.410 41.450 61.910 41.620 ;
        RECT 62.790 41.450 63.290 41.620 ;
        RECT 64.170 41.450 64.670 41.620 ;
        RECT 65.550 41.450 66.050 41.620 ;
        RECT 66.930 41.450 67.430 41.620 ;
        RECT 68.310 41.450 68.810 41.620 ;
        RECT 55.890 40.910 56.390 41.080 ;
        RECT 57.270 40.910 57.770 41.080 ;
        RECT 58.650 40.910 59.150 41.080 ;
        RECT 60.030 40.910 60.530 41.080 ;
        RECT 61.410 40.910 61.910 41.080 ;
        RECT 62.790 40.910 63.290 41.080 ;
        RECT 64.170 40.910 64.670 41.080 ;
        RECT 65.550 40.910 66.050 41.080 ;
        RECT 66.930 40.910 67.430 41.080 ;
        RECT 68.310 40.910 68.810 41.080 ;
        RECT 55.660 40.050 55.830 40.740 ;
        RECT 56.450 40.050 56.620 40.740 ;
        RECT 57.040 40.050 57.210 40.740 ;
        RECT 57.830 40.050 58.000 40.740 ;
        RECT 58.420 40.050 58.590 40.740 ;
        RECT 59.210 40.050 59.380 40.740 ;
        RECT 59.800 40.050 59.970 40.740 ;
        RECT 60.590 40.050 60.760 40.740 ;
        RECT 61.180 40.050 61.350 40.740 ;
        RECT 61.970 40.050 62.140 40.740 ;
        RECT 62.560 40.050 62.730 40.740 ;
        RECT 63.350 40.050 63.520 40.740 ;
        RECT 63.940 40.050 64.110 40.740 ;
        RECT 64.730 40.050 64.900 40.740 ;
        RECT 65.320 40.050 65.490 40.740 ;
        RECT 66.110 40.050 66.280 40.740 ;
        RECT 66.700 40.050 66.870 40.740 ;
        RECT 67.490 40.050 67.660 40.740 ;
        RECT 68.080 40.050 68.250 40.740 ;
        RECT 68.870 40.050 69.040 40.740 ;
        RECT 55.890 39.710 56.390 39.880 ;
        RECT 57.270 39.710 57.770 39.880 ;
        RECT 58.650 39.710 59.150 39.880 ;
        RECT 60.030 39.710 60.530 39.880 ;
        RECT 61.410 39.710 61.910 39.880 ;
        RECT 62.790 39.710 63.290 39.880 ;
        RECT 64.170 39.710 64.670 39.880 ;
        RECT 65.550 39.710 66.050 39.880 ;
        RECT 66.930 39.710 67.430 39.880 ;
        RECT 68.310 39.710 68.810 39.880 ;
        RECT 69.530 39.415 69.700 43.115 ;
        RECT 54.950 39.245 69.700 39.415 ;
        RECT 55.980 37.910 56.980 38.080 ;
        RECT 57.290 38.015 57.500 38.385 ;
        RECT 57.860 37.910 58.860 38.080 ;
        RECT 59.170 38.015 59.380 38.385 ;
        RECT 59.740 37.910 60.740 38.080 ;
        RECT 61.050 38.015 61.260 38.385 ;
        RECT 61.620 37.910 62.620 38.080 ;
        RECT 62.930 38.015 63.140 38.385 ;
        RECT 63.500 37.910 64.500 38.080 ;
        RECT 64.810 38.015 65.020 38.385 ;
        RECT 65.380 37.910 66.380 38.080 ;
        RECT 33.120 37.710 47.320 37.880 ;
        RECT 33.020 36.660 47.470 36.830 ;
        RECT 33.020 34.700 33.190 36.660 ;
        RECT 33.970 36.195 34.470 36.365 ;
        RECT 35.470 36.195 35.970 36.365 ;
        RECT 36.970 36.195 37.470 36.365 ;
        RECT 38.470 36.195 38.970 36.365 ;
        RECT 39.970 36.195 40.470 36.365 ;
        RECT 41.470 36.195 41.970 36.365 ;
        RECT 42.970 36.195 43.470 36.365 ;
        RECT 44.470 36.195 44.970 36.365 ;
        RECT 45.970 36.195 46.470 36.365 ;
        RECT 33.680 35.335 33.850 36.025 ;
        RECT 34.590 35.335 34.760 36.025 ;
        RECT 35.180 35.335 35.350 36.025 ;
        RECT 36.090 35.335 36.260 36.025 ;
        RECT 36.680 35.335 36.850 36.025 ;
        RECT 37.590 35.335 37.760 36.025 ;
        RECT 38.180 35.335 38.350 36.025 ;
        RECT 39.090 35.335 39.260 36.025 ;
        RECT 39.680 35.335 39.850 36.025 ;
        RECT 40.590 35.335 40.760 36.025 ;
        RECT 41.180 35.335 41.350 36.025 ;
        RECT 42.090 35.335 42.260 36.025 ;
        RECT 42.680 35.335 42.850 36.025 ;
        RECT 43.590 35.335 43.760 36.025 ;
        RECT 44.180 35.335 44.350 36.025 ;
        RECT 45.090 35.335 45.260 36.025 ;
        RECT 45.680 35.335 45.850 36.025 ;
        RECT 46.590 35.335 46.760 36.025 ;
        RECT 33.970 34.995 34.470 35.165 ;
        RECT 35.470 34.995 35.970 35.165 ;
        RECT 36.970 34.995 37.470 35.165 ;
        RECT 38.470 34.995 38.970 35.165 ;
        RECT 39.970 34.995 40.470 35.165 ;
        RECT 41.470 34.995 41.970 35.165 ;
        RECT 42.970 34.995 43.470 35.165 ;
        RECT 44.470 34.995 44.970 35.165 ;
        RECT 45.970 34.995 46.470 35.165 ;
        RECT 47.300 34.700 47.470 36.660 ;
        RECT 33.020 34.530 47.470 34.700 ;
        RECT 55.750 33.655 55.920 37.695 ;
        RECT 57.040 33.655 57.210 37.695 ;
        RECT 57.630 33.655 57.800 37.695 ;
        RECT 58.920 33.655 59.090 37.695 ;
        RECT 59.510 33.655 59.680 37.695 ;
        RECT 60.800 33.655 60.970 37.695 ;
        RECT 61.390 33.655 61.560 37.695 ;
        RECT 62.680 33.655 62.850 37.695 ;
        RECT 63.270 33.655 63.440 37.695 ;
        RECT 64.560 33.655 64.730 37.695 ;
        RECT 65.150 33.655 65.320 37.695 ;
        RECT 66.440 33.655 66.610 37.695 ;
        RECT 67.150 36.515 67.500 38.675 ;
        RECT 67.980 36.515 68.330 38.675 ;
        RECT 68.810 36.515 69.160 38.675 ;
        RECT 69.640 36.515 69.990 38.675 ;
        RECT 55.980 33.270 56.980 33.440 ;
        RECT 57.860 33.270 58.860 33.440 ;
        RECT 59.740 33.270 60.740 33.440 ;
        RECT 61.620 33.270 62.620 33.440 ;
        RECT 63.500 33.270 64.500 33.440 ;
        RECT 65.380 33.270 66.380 33.440 ;
        RECT 55.980 32.730 56.980 32.900 ;
        RECT 57.860 32.730 58.860 32.900 ;
        RECT 59.740 32.730 60.740 32.900 ;
        RECT 61.620 32.730 62.620 32.900 ;
        RECT 63.500 32.730 64.500 32.900 ;
        RECT 65.380 32.730 66.380 32.900 ;
        RECT 55.750 28.475 55.920 32.515 ;
        RECT 57.040 28.475 57.210 32.515 ;
        RECT 57.630 28.475 57.800 32.515 ;
        RECT 58.920 28.475 59.090 32.515 ;
        RECT 59.510 28.475 59.680 32.515 ;
        RECT 60.800 28.475 60.970 32.515 ;
        RECT 61.390 28.475 61.560 32.515 ;
        RECT 62.680 28.475 62.850 32.515 ;
        RECT 63.270 28.475 63.440 32.515 ;
        RECT 64.560 28.475 64.730 32.515 ;
        RECT 65.150 28.475 65.320 32.515 ;
        RECT 66.440 28.475 66.610 32.515 ;
        RECT 67.150 28.265 67.500 30.425 ;
        RECT 67.980 28.265 68.330 30.425 ;
        RECT 68.810 28.265 69.160 30.425 ;
        RECT 69.640 28.265 69.990 30.425 ;
        RECT 55.980 28.090 56.980 28.260 ;
        RECT 57.860 28.090 58.860 28.260 ;
        RECT 59.740 28.090 60.740 28.260 ;
        RECT 61.620 28.090 62.620 28.260 ;
        RECT 63.500 28.090 64.500 28.260 ;
        RECT 65.380 28.090 66.380 28.260 ;
        RECT 55.980 27.535 56.980 27.705 ;
        RECT 57.860 27.535 58.860 27.705 ;
        RECT 59.740 27.535 60.740 27.705 ;
        RECT 61.620 27.535 62.620 27.705 ;
        RECT 63.500 27.535 64.500 27.705 ;
        RECT 65.380 27.535 66.380 27.705 ;
        RECT 67.260 27.535 68.260 27.705 ;
        RECT 55.750 25.325 55.920 27.365 ;
        RECT 57.040 25.325 57.210 27.365 ;
        RECT 57.630 25.325 57.800 27.365 ;
        RECT 58.920 25.325 59.090 27.365 ;
        RECT 59.510 25.325 59.680 27.365 ;
        RECT 60.800 25.325 60.970 27.365 ;
        RECT 61.390 25.325 61.560 27.365 ;
        RECT 62.680 25.325 62.850 27.365 ;
        RECT 63.270 25.325 63.440 27.365 ;
        RECT 64.560 25.325 64.730 27.365 ;
        RECT 65.150 25.325 65.320 27.365 ;
        RECT 66.440 25.325 66.610 27.365 ;
        RECT 67.030 25.325 67.200 27.365 ;
        RECT 68.320 25.325 68.490 27.365 ;
        RECT 69.750 26.585 69.960 26.955 ;
        RECT 69.750 25.300 69.960 25.670 ;
        RECT 55.980 24.985 56.980 25.155 ;
        RECT 57.860 24.985 58.860 25.155 ;
        RECT 59.740 24.985 60.740 25.155 ;
        RECT 61.620 24.985 62.620 25.155 ;
        RECT 63.500 24.985 64.500 25.155 ;
        RECT 65.380 24.985 66.380 25.155 ;
        RECT 67.260 24.985 68.260 25.155 ;
        RECT 55.980 24.445 56.980 24.615 ;
        RECT 57.860 24.445 58.860 24.615 ;
        RECT 59.740 24.445 60.740 24.615 ;
        RECT 61.620 24.445 62.620 24.615 ;
        RECT 63.500 24.445 64.500 24.615 ;
        RECT 65.380 24.445 66.380 24.615 ;
        RECT 67.260 24.445 68.260 24.615 ;
        RECT 55.750 22.235 55.920 24.275 ;
        RECT 57.040 22.235 57.210 24.275 ;
        RECT 57.630 22.235 57.800 24.275 ;
        RECT 58.920 22.235 59.090 24.275 ;
        RECT 59.510 22.235 59.680 24.275 ;
        RECT 60.800 22.235 60.970 24.275 ;
        RECT 61.390 22.235 61.560 24.275 ;
        RECT 62.680 22.235 62.850 24.275 ;
        RECT 63.270 22.235 63.440 24.275 ;
        RECT 64.560 22.235 64.730 24.275 ;
        RECT 65.150 22.235 65.320 24.275 ;
        RECT 66.440 22.235 66.610 24.275 ;
        RECT 67.030 22.235 67.200 24.275 ;
        RECT 68.320 22.235 68.490 24.275 ;
        RECT 69.750 24.015 69.960 24.385 ;
        RECT 69.750 22.725 69.960 23.095 ;
        RECT 55.980 21.895 56.980 22.065 ;
        RECT 57.860 21.895 58.860 22.065 ;
        RECT 59.740 21.895 60.740 22.065 ;
        RECT 61.620 21.895 62.620 22.065 ;
        RECT 63.500 21.895 64.500 22.065 ;
        RECT 65.380 21.895 66.380 22.065 ;
        RECT 67.260 21.895 68.260 22.065 ;
        RECT 72.965 20.455 73.135 104.115 ;
        RECT 99.920 75.735 122.720 75.905 ;
        RECT 29.585 20.285 73.135 20.455 ;
        RECT 82.285 35.430 91.435 35.600 ;
        RECT 82.285 20.455 82.455 35.430 ;
        RECT 85.820 31.895 87.900 32.065 ;
        RECT 85.820 27.405 85.990 31.895 ;
        RECT 86.610 31.475 87.110 31.645 ;
        RECT 86.380 30.220 86.550 31.260 ;
        RECT 87.170 30.220 87.340 31.260 ;
        RECT 86.610 29.835 87.110 30.005 ;
        RECT 86.610 29.295 87.110 29.465 ;
        RECT 86.380 28.040 86.550 29.080 ;
        RECT 87.170 28.040 87.340 29.080 ;
        RECT 86.610 27.655 87.110 27.825 ;
        RECT 87.730 27.405 87.900 31.895 ;
        RECT 85.820 27.235 87.900 27.405 ;
        RECT 85.720 26.185 88.050 26.355 ;
        RECT 85.720 22.485 85.890 26.185 ;
        RECT 86.610 25.720 87.110 25.890 ;
        RECT 86.380 24.860 86.550 25.550 ;
        RECT 87.170 24.860 87.340 25.550 ;
        RECT 86.610 24.520 87.110 24.690 ;
        RECT 86.610 23.980 87.110 24.150 ;
        RECT 86.380 23.120 86.550 23.810 ;
        RECT 87.170 23.120 87.340 23.810 ;
        RECT 86.610 22.780 87.110 22.950 ;
        RECT 87.880 22.485 88.050 26.185 ;
        RECT 85.720 22.315 88.050 22.485 ;
        RECT 91.265 20.455 91.435 35.430 ;
        RECT 82.285 20.285 91.435 20.455 ;
        RECT 99.920 20.455 100.090 75.735 ;
        RECT 102.225 72.950 102.575 75.110 ;
        RECT 103.055 72.950 103.405 75.110 ;
        RECT 103.885 72.950 104.235 75.110 ;
        RECT 104.715 72.950 105.065 75.110 ;
        RECT 105.545 72.950 105.895 75.110 ;
        RECT 106.375 72.950 106.725 75.110 ;
        RECT 107.205 72.950 107.555 75.110 ;
        RECT 108.035 72.950 108.385 75.110 ;
        RECT 108.865 72.950 109.215 75.110 ;
        RECT 109.695 72.950 110.045 75.110 ;
        RECT 110.525 72.950 110.875 75.110 ;
        RECT 111.355 72.950 111.705 75.110 ;
        RECT 112.185 72.950 112.535 75.110 ;
        RECT 113.015 72.950 113.365 75.110 ;
        RECT 113.845 72.950 114.195 75.110 ;
        RECT 114.675 72.950 115.025 75.110 ;
        RECT 115.505 72.950 115.855 75.110 ;
        RECT 116.335 72.950 116.685 75.110 ;
        RECT 117.165 72.950 117.515 75.110 ;
        RECT 117.995 72.950 118.345 75.110 ;
        RECT 118.825 72.950 119.175 75.110 ;
        RECT 119.655 72.950 120.005 75.110 ;
        RECT 120.485 72.950 120.835 75.110 ;
        RECT 121.315 72.950 121.665 75.110 ;
        RECT 102.225 38.950 102.575 41.110 ;
        RECT 103.055 38.950 103.405 41.110 ;
        RECT 103.885 38.950 104.235 41.110 ;
        RECT 104.715 38.950 105.065 41.110 ;
        RECT 105.545 38.950 105.895 41.110 ;
        RECT 106.375 38.950 106.725 41.110 ;
        RECT 107.205 38.950 107.555 41.110 ;
        RECT 108.035 38.950 108.385 41.110 ;
        RECT 108.865 38.950 109.215 41.110 ;
        RECT 109.695 38.950 110.045 41.110 ;
        RECT 110.525 38.950 110.875 41.110 ;
        RECT 111.355 38.950 111.705 41.110 ;
        RECT 112.185 38.950 112.535 41.110 ;
        RECT 113.015 38.950 113.365 41.110 ;
        RECT 113.845 38.950 114.195 41.110 ;
        RECT 114.675 38.950 115.025 41.110 ;
        RECT 115.505 38.950 115.855 41.110 ;
        RECT 116.335 38.950 116.685 41.110 ;
        RECT 117.165 38.950 117.515 41.110 ;
        RECT 117.995 38.950 118.345 41.110 ;
        RECT 118.825 38.950 119.175 41.110 ;
        RECT 119.655 38.950 120.005 41.110 ;
        RECT 120.485 38.950 120.835 41.110 ;
        RECT 121.315 38.950 121.665 41.110 ;
        RECT 102.225 36.515 102.575 38.675 ;
        RECT 103.055 36.515 103.405 38.675 ;
        RECT 103.885 36.515 104.235 38.675 ;
        RECT 104.715 36.515 105.065 38.675 ;
        RECT 105.835 37.910 106.835 38.080 ;
        RECT 107.195 38.015 107.405 38.385 ;
        RECT 107.715 37.910 108.715 38.080 ;
        RECT 109.075 38.015 109.285 38.385 ;
        RECT 109.595 37.910 110.595 38.080 ;
        RECT 110.955 38.015 111.165 38.385 ;
        RECT 111.475 37.910 112.475 38.080 ;
        RECT 112.835 38.015 113.045 38.385 ;
        RECT 113.355 37.910 114.355 38.080 ;
        RECT 114.715 38.015 114.925 38.385 ;
        RECT 115.235 37.910 116.235 38.080 ;
        RECT 105.605 33.655 105.775 37.695 ;
        RECT 106.895 33.655 107.065 37.695 ;
        RECT 107.485 33.655 107.655 37.695 ;
        RECT 108.775 33.655 108.945 37.695 ;
        RECT 109.365 33.655 109.535 37.695 ;
        RECT 110.655 33.655 110.825 37.695 ;
        RECT 111.245 33.655 111.415 37.695 ;
        RECT 112.535 33.655 112.705 37.695 ;
        RECT 113.125 33.655 113.295 37.695 ;
        RECT 114.415 33.655 114.585 37.695 ;
        RECT 115.005 33.655 115.175 37.695 ;
        RECT 116.295 33.655 116.465 37.695 ;
        RECT 105.835 33.270 106.835 33.440 ;
        RECT 107.715 33.270 108.715 33.440 ;
        RECT 109.595 33.270 110.595 33.440 ;
        RECT 111.475 33.270 112.475 33.440 ;
        RECT 113.355 33.270 114.355 33.440 ;
        RECT 115.235 33.270 116.235 33.440 ;
        RECT 105.835 32.730 106.835 32.900 ;
        RECT 107.715 32.730 108.715 32.900 ;
        RECT 109.595 32.730 110.595 32.900 ;
        RECT 111.475 32.730 112.475 32.900 ;
        RECT 113.355 32.730 114.355 32.900 ;
        RECT 115.235 32.730 116.235 32.900 ;
        RECT 102.225 28.265 102.575 30.425 ;
        RECT 103.055 28.265 103.405 30.425 ;
        RECT 103.885 28.265 104.235 30.425 ;
        RECT 104.715 28.265 105.065 30.425 ;
        RECT 105.605 28.475 105.775 32.515 ;
        RECT 106.895 28.475 107.065 32.515 ;
        RECT 107.485 28.475 107.655 32.515 ;
        RECT 108.775 28.475 108.945 32.515 ;
        RECT 109.365 28.475 109.535 32.515 ;
        RECT 110.655 28.475 110.825 32.515 ;
        RECT 111.245 28.475 111.415 32.515 ;
        RECT 112.535 28.475 112.705 32.515 ;
        RECT 113.125 28.475 113.295 32.515 ;
        RECT 114.415 28.475 114.585 32.515 ;
        RECT 115.005 28.475 115.175 32.515 ;
        RECT 116.295 28.475 116.465 32.515 ;
        RECT 105.835 28.090 106.835 28.260 ;
        RECT 107.715 28.090 108.715 28.260 ;
        RECT 109.595 28.090 110.595 28.260 ;
        RECT 111.475 28.090 112.475 28.260 ;
        RECT 113.355 28.090 114.355 28.260 ;
        RECT 115.235 28.090 116.235 28.260 ;
        RECT 103.955 27.535 104.955 27.705 ;
        RECT 105.835 27.535 106.835 27.705 ;
        RECT 107.715 27.535 108.715 27.705 ;
        RECT 109.595 27.535 110.595 27.705 ;
        RECT 111.475 27.535 112.475 27.705 ;
        RECT 113.355 27.535 114.355 27.705 ;
        RECT 115.235 27.535 116.235 27.705 ;
        RECT 102.255 26.585 102.465 26.955 ;
        RECT 102.255 25.300 102.465 25.670 ;
        RECT 103.725 25.325 103.895 27.365 ;
        RECT 105.015 25.325 105.185 27.365 ;
        RECT 105.605 25.325 105.775 27.365 ;
        RECT 106.895 25.325 107.065 27.365 ;
        RECT 107.485 25.325 107.655 27.365 ;
        RECT 108.775 25.325 108.945 27.365 ;
        RECT 109.365 25.325 109.535 27.365 ;
        RECT 110.655 25.325 110.825 27.365 ;
        RECT 111.245 25.325 111.415 27.365 ;
        RECT 112.535 25.325 112.705 27.365 ;
        RECT 113.125 25.325 113.295 27.365 ;
        RECT 114.415 25.325 114.585 27.365 ;
        RECT 115.005 25.325 115.175 27.365 ;
        RECT 116.295 25.325 116.465 27.365 ;
        RECT 103.955 24.985 104.955 25.155 ;
        RECT 105.835 24.985 106.835 25.155 ;
        RECT 107.715 24.985 108.715 25.155 ;
        RECT 109.595 24.985 110.595 25.155 ;
        RECT 111.475 24.985 112.475 25.155 ;
        RECT 113.355 24.985 114.355 25.155 ;
        RECT 115.235 24.985 116.235 25.155 ;
        RECT 103.955 24.445 104.955 24.615 ;
        RECT 105.835 24.445 106.835 24.615 ;
        RECT 107.715 24.445 108.715 24.615 ;
        RECT 109.595 24.445 110.595 24.615 ;
        RECT 111.475 24.445 112.475 24.615 ;
        RECT 113.355 24.445 114.355 24.615 ;
        RECT 115.235 24.445 116.235 24.615 ;
        RECT 102.255 24.015 102.465 24.385 ;
        RECT 102.255 22.725 102.465 23.095 ;
        RECT 103.725 22.235 103.895 24.275 ;
        RECT 105.015 22.235 105.185 24.275 ;
        RECT 105.605 22.235 105.775 24.275 ;
        RECT 106.895 22.235 107.065 24.275 ;
        RECT 107.485 22.235 107.655 24.275 ;
        RECT 108.775 22.235 108.945 24.275 ;
        RECT 109.365 22.235 109.535 24.275 ;
        RECT 110.655 22.235 110.825 24.275 ;
        RECT 111.245 22.235 111.415 24.275 ;
        RECT 112.535 22.235 112.705 24.275 ;
        RECT 113.125 22.235 113.295 24.275 ;
        RECT 114.415 22.235 114.585 24.275 ;
        RECT 115.005 22.235 115.175 24.275 ;
        RECT 116.295 22.235 116.465 24.275 ;
        RECT 103.955 21.895 104.955 22.065 ;
        RECT 105.835 21.895 106.835 22.065 ;
        RECT 107.715 21.895 108.715 22.065 ;
        RECT 109.595 21.895 110.595 22.065 ;
        RECT 111.475 21.895 112.475 22.065 ;
        RECT 113.355 21.895 114.355 22.065 ;
        RECT 115.235 21.895 116.235 22.065 ;
        RECT 122.550 20.455 122.720 75.735 ;
        RECT 99.920 20.285 122.720 20.455 ;
      LAYER met1 ;
        RECT 0.000 224.760 1.000 225.760 ;
        RECT 144.360 224.760 145.360 225.760 ;
        RECT 38.610 208.130 38.900 208.160 ;
        RECT 40.250 208.130 40.510 208.145 ;
        RECT 41.750 208.130 42.010 208.145 ;
        RECT 43.250 208.130 43.510 208.145 ;
        RECT 44.750 208.130 45.010 208.145 ;
        RECT 46.250 208.130 46.510 208.145 ;
        RECT 47.750 208.130 48.010 208.145 ;
        RECT 49.250 208.130 49.510 208.145 ;
        RECT 50.750 208.130 51.010 208.145 ;
        RECT 51.390 208.130 51.680 208.160 ;
        RECT 38.610 207.840 51.680 208.130 ;
        RECT 38.610 207.810 38.900 207.840 ;
        RECT 40.250 207.825 40.510 207.840 ;
        RECT 41.750 207.825 42.010 207.840 ;
        RECT 43.250 207.825 43.510 207.840 ;
        RECT 44.750 207.825 45.010 207.840 ;
        RECT 46.250 207.825 46.510 207.840 ;
        RECT 47.750 207.825 48.010 207.840 ;
        RECT 49.250 207.825 49.510 207.840 ;
        RECT 50.750 207.825 51.010 207.840 ;
        RECT 39.690 207.405 40.150 207.635 ;
        RECT 39.380 207.260 39.550 207.265 ;
        RECT 39.335 207.230 39.595 207.260 ;
        RECT 39.305 206.970 39.625 207.230 ;
        RECT 39.335 206.940 39.595 206.970 ;
        RECT 13.320 206.705 13.620 206.740 ;
        RECT 14.820 206.705 15.120 206.740 ;
        RECT 16.320 206.705 16.620 206.740 ;
        RECT 17.820 206.705 18.120 206.740 ;
        RECT 19.320 206.705 19.620 206.740 ;
        RECT 20.820 206.705 21.120 206.740 ;
        RECT 22.320 206.705 22.620 206.740 ;
        RECT 23.820 206.705 24.120 206.740 ;
        RECT 13.170 206.415 25.170 206.705 ;
        RECT 39.350 206.595 39.580 206.940 ;
        RECT 13.320 206.380 13.620 206.415 ;
        RECT 14.820 206.380 15.120 206.415 ;
        RECT 16.320 206.380 16.620 206.415 ;
        RECT 17.820 206.380 18.120 206.415 ;
        RECT 19.320 206.380 19.620 206.415 ;
        RECT 20.820 206.380 21.120 206.415 ;
        RECT 22.320 206.380 22.620 206.415 ;
        RECT 23.820 206.380 24.120 206.415 ;
        RECT 13.380 205.820 13.550 206.380 ;
        RECT 13.690 206.025 14.150 206.255 ;
        RECT 13.350 204.820 13.580 205.820 ;
        RECT 13.380 204.800 13.550 204.820 ;
        RECT 13.835 204.615 14.005 206.025 ;
        RECT 14.170 205.500 14.580 205.850 ;
        RECT 14.880 205.820 15.050 206.380 ;
        RECT 15.190 206.025 15.650 206.255 ;
        RECT 14.260 204.820 14.490 205.500 ;
        RECT 14.850 204.820 15.080 205.820 ;
        RECT 14.290 204.800 14.460 204.820 ;
        RECT 14.880 204.800 15.050 204.820 ;
        RECT 15.335 204.615 15.505 206.025 ;
        RECT 15.670 205.500 16.080 205.850 ;
        RECT 16.380 205.820 16.550 206.380 ;
        RECT 16.690 206.025 17.150 206.255 ;
        RECT 15.760 204.820 15.990 205.500 ;
        RECT 16.350 204.820 16.580 205.820 ;
        RECT 15.790 204.800 15.960 204.820 ;
        RECT 16.380 204.800 16.550 204.820 ;
        RECT 16.835 204.615 17.005 206.025 ;
        RECT 17.170 205.500 17.580 205.850 ;
        RECT 17.880 205.820 18.050 206.380 ;
        RECT 18.190 206.025 18.650 206.255 ;
        RECT 17.260 204.820 17.490 205.500 ;
        RECT 17.850 204.820 18.080 205.820 ;
        RECT 17.290 204.800 17.460 204.820 ;
        RECT 17.880 204.800 18.050 204.820 ;
        RECT 18.335 204.615 18.505 206.025 ;
        RECT 18.670 205.500 19.080 205.850 ;
        RECT 19.380 205.820 19.550 206.380 ;
        RECT 19.690 206.025 20.150 206.255 ;
        RECT 18.760 204.820 18.990 205.500 ;
        RECT 19.350 204.820 19.580 205.820 ;
        RECT 18.790 204.800 18.960 204.820 ;
        RECT 19.380 204.800 19.550 204.820 ;
        RECT 19.835 204.615 20.005 206.025 ;
        RECT 20.170 205.500 20.580 205.850 ;
        RECT 20.880 205.820 21.050 206.380 ;
        RECT 21.190 206.025 21.650 206.255 ;
        RECT 20.260 204.820 20.490 205.500 ;
        RECT 20.850 204.820 21.080 205.820 ;
        RECT 20.290 204.800 20.460 204.820 ;
        RECT 20.880 204.800 21.050 204.820 ;
        RECT 21.335 204.615 21.505 206.025 ;
        RECT 21.670 205.500 22.080 205.850 ;
        RECT 22.380 205.820 22.550 206.380 ;
        RECT 22.690 206.025 23.150 206.255 ;
        RECT 21.760 204.820 21.990 205.500 ;
        RECT 22.350 204.820 22.580 205.820 ;
        RECT 21.790 204.800 21.960 204.820 ;
        RECT 22.380 204.800 22.550 204.820 ;
        RECT 22.835 204.615 23.005 206.025 ;
        RECT 23.170 205.500 23.580 205.850 ;
        RECT 23.880 205.820 24.050 206.380 ;
        RECT 24.190 206.025 24.650 206.255 ;
        RECT 23.260 204.820 23.490 205.500 ;
        RECT 23.850 204.820 24.080 205.820 ;
        RECT 23.290 204.800 23.460 204.820 ;
        RECT 23.880 204.800 24.050 204.820 ;
        RECT 24.335 204.615 24.505 206.025 ;
        RECT 24.670 205.500 25.080 205.850 ;
        RECT 24.760 204.820 24.990 205.500 ;
        RECT 24.790 204.800 24.960 204.820 ;
        RECT 13.690 204.385 14.150 204.615 ;
        RECT 15.190 204.385 15.650 204.615 ;
        RECT 16.690 204.385 17.150 204.615 ;
        RECT 18.190 204.385 18.650 204.615 ;
        RECT 19.690 204.385 20.150 204.615 ;
        RECT 21.190 204.385 21.650 204.615 ;
        RECT 22.690 204.385 23.150 204.615 ;
        RECT 24.190 204.385 24.650 204.615 ;
        RECT 13.835 202.680 14.005 204.385 ;
        RECT 15.335 202.680 15.505 204.385 ;
        RECT 16.835 202.680 17.005 204.385 ;
        RECT 18.335 202.680 18.505 204.385 ;
        RECT 19.835 202.680 20.005 204.385 ;
        RECT 21.335 202.680 21.505 204.385 ;
        RECT 22.835 202.680 23.005 204.385 ;
        RECT 24.335 202.680 24.505 204.385 ;
        RECT 39.380 204.065 39.550 206.595 ;
        RECT 39.835 206.480 40.005 207.405 ;
        RECT 40.290 207.245 40.460 207.825 ;
        RECT 41.190 207.405 41.650 207.635 ;
        RECT 40.880 207.260 41.050 207.265 ;
        RECT 40.260 206.595 40.490 207.245 ;
        RECT 40.835 207.230 41.095 207.260 ;
        RECT 40.805 206.970 41.125 207.230 ;
        RECT 40.835 206.940 41.095 206.970 ;
        RECT 40.850 206.595 41.080 206.940 ;
        RECT 40.290 206.575 40.460 206.595 ;
        RECT 39.790 206.435 40.050 206.480 ;
        RECT 39.690 206.205 40.150 206.435 ;
        RECT 39.790 206.160 40.050 206.205 ;
        RECT 39.690 204.270 40.150 204.500 ;
        RECT 39.350 203.360 39.580 204.065 ;
        RECT 39.305 203.100 39.625 203.360 ;
        RECT 39.350 203.065 39.580 203.100 ;
        RECT 39.380 203.045 39.550 203.065 ;
        RECT 39.210 202.830 39.530 202.875 ;
        RECT 39.835 202.860 40.005 204.270 ;
        RECT 40.290 204.065 40.460 204.085 ;
        RECT 40.880 204.065 41.050 206.595 ;
        RECT 41.335 206.480 41.505 207.405 ;
        RECT 41.790 207.245 41.960 207.825 ;
        RECT 42.690 207.405 43.150 207.635 ;
        RECT 42.380 207.260 42.550 207.265 ;
        RECT 41.760 206.595 41.990 207.245 ;
        RECT 42.335 207.230 42.595 207.260 ;
        RECT 42.305 206.970 42.625 207.230 ;
        RECT 42.335 206.940 42.595 206.970 ;
        RECT 42.350 206.595 42.580 206.940 ;
        RECT 41.790 206.575 41.960 206.595 ;
        RECT 41.290 206.435 41.550 206.480 ;
        RECT 41.190 206.205 41.650 206.435 ;
        RECT 41.290 206.160 41.550 206.205 ;
        RECT 41.190 204.270 41.650 204.500 ;
        RECT 40.260 203.065 40.490 204.065 ;
        RECT 40.850 203.360 41.080 204.065 ;
        RECT 40.805 203.100 41.125 203.360 ;
        RECT 40.850 203.065 41.080 203.100 ;
        RECT 39.690 202.830 40.150 202.860 ;
        RECT 13.690 202.450 14.150 202.680 ;
        RECT 15.190 202.450 15.650 202.680 ;
        RECT 16.690 202.450 17.150 202.680 ;
        RECT 18.190 202.450 18.650 202.680 ;
        RECT 19.690 202.450 20.150 202.680 ;
        RECT 21.190 202.450 21.650 202.680 ;
        RECT 22.690 202.450 23.150 202.680 ;
        RECT 24.190 202.450 24.650 202.680 ;
        RECT 39.210 202.660 40.150 202.830 ;
        RECT 39.210 202.615 39.530 202.660 ;
        RECT 39.690 202.630 40.150 202.660 ;
        RECT 38.725 202.470 39.075 202.530 ;
        RECT 40.290 202.470 40.460 203.065 ;
        RECT 40.880 203.045 41.050 203.065 ;
        RECT 40.710 202.830 41.030 202.875 ;
        RECT 41.335 202.860 41.505 204.270 ;
        RECT 41.790 204.065 41.960 204.085 ;
        RECT 42.380 204.065 42.550 206.595 ;
        RECT 42.835 206.480 43.005 207.405 ;
        RECT 43.290 207.245 43.460 207.825 ;
        RECT 44.190 207.405 44.650 207.635 ;
        RECT 43.880 207.260 44.050 207.265 ;
        RECT 43.260 206.595 43.490 207.245 ;
        RECT 43.835 207.230 44.095 207.260 ;
        RECT 43.805 206.970 44.125 207.230 ;
        RECT 43.835 206.940 44.095 206.970 ;
        RECT 43.850 206.595 44.080 206.940 ;
        RECT 43.290 206.575 43.460 206.595 ;
        RECT 42.790 206.435 43.050 206.480 ;
        RECT 42.690 206.205 43.150 206.435 ;
        RECT 42.790 206.160 43.050 206.205 ;
        RECT 42.690 204.270 43.150 204.500 ;
        RECT 41.760 203.065 41.990 204.065 ;
        RECT 42.350 203.360 42.580 204.065 ;
        RECT 42.305 203.100 42.625 203.360 ;
        RECT 42.350 203.065 42.580 203.100 ;
        RECT 41.190 202.830 41.650 202.860 ;
        RECT 40.710 202.660 41.650 202.830 ;
        RECT 40.710 202.615 41.030 202.660 ;
        RECT 41.190 202.630 41.650 202.660 ;
        RECT 41.790 202.470 41.960 203.065 ;
        RECT 42.380 203.045 42.550 203.065 ;
        RECT 42.210 202.830 42.530 202.875 ;
        RECT 42.835 202.860 43.005 204.270 ;
        RECT 43.290 204.065 43.460 204.085 ;
        RECT 43.880 204.065 44.050 206.595 ;
        RECT 44.335 206.480 44.505 207.405 ;
        RECT 44.790 207.245 44.960 207.825 ;
        RECT 45.690 207.405 46.150 207.635 ;
        RECT 45.380 207.260 45.550 207.265 ;
        RECT 44.760 206.595 44.990 207.245 ;
        RECT 45.335 207.230 45.595 207.260 ;
        RECT 45.305 206.970 45.625 207.230 ;
        RECT 45.335 206.940 45.595 206.970 ;
        RECT 45.350 206.595 45.580 206.940 ;
        RECT 44.790 206.575 44.960 206.595 ;
        RECT 44.290 206.435 44.550 206.480 ;
        RECT 44.190 206.205 44.650 206.435 ;
        RECT 44.290 206.160 44.550 206.205 ;
        RECT 44.190 204.270 44.650 204.500 ;
        RECT 43.260 203.065 43.490 204.065 ;
        RECT 43.850 203.360 44.080 204.065 ;
        RECT 43.805 203.100 44.125 203.360 ;
        RECT 43.850 203.065 44.080 203.100 ;
        RECT 42.690 202.830 43.150 202.860 ;
        RECT 42.210 202.660 43.150 202.830 ;
        RECT 42.210 202.615 42.530 202.660 ;
        RECT 42.690 202.630 43.150 202.660 ;
        RECT 43.290 202.470 43.460 203.065 ;
        RECT 43.880 203.045 44.050 203.065 ;
        RECT 43.710 202.830 44.030 202.875 ;
        RECT 44.335 202.860 44.505 204.270 ;
        RECT 44.790 204.065 44.960 204.085 ;
        RECT 45.380 204.065 45.550 206.595 ;
        RECT 45.835 206.480 46.005 207.405 ;
        RECT 46.290 207.245 46.460 207.825 ;
        RECT 47.190 207.405 47.650 207.635 ;
        RECT 46.880 207.260 47.050 207.265 ;
        RECT 46.260 206.595 46.490 207.245 ;
        RECT 46.835 207.230 47.095 207.260 ;
        RECT 46.805 206.970 47.125 207.230 ;
        RECT 46.835 206.940 47.095 206.970 ;
        RECT 46.850 206.595 47.080 206.940 ;
        RECT 46.290 206.575 46.460 206.595 ;
        RECT 45.790 206.435 46.050 206.480 ;
        RECT 45.690 206.205 46.150 206.435 ;
        RECT 45.790 206.160 46.050 206.205 ;
        RECT 45.690 204.270 46.150 204.500 ;
        RECT 44.760 203.065 44.990 204.065 ;
        RECT 45.350 203.360 45.580 204.065 ;
        RECT 45.305 203.100 45.625 203.360 ;
        RECT 45.350 203.065 45.580 203.100 ;
        RECT 44.190 202.830 44.650 202.860 ;
        RECT 43.710 202.660 44.650 202.830 ;
        RECT 43.710 202.615 44.030 202.660 ;
        RECT 44.190 202.630 44.650 202.660 ;
        RECT 44.790 202.470 44.960 203.065 ;
        RECT 45.380 203.045 45.550 203.065 ;
        RECT 45.210 202.830 45.530 202.875 ;
        RECT 45.835 202.860 46.005 204.270 ;
        RECT 46.290 204.065 46.460 204.085 ;
        RECT 46.880 204.065 47.050 206.595 ;
        RECT 47.335 206.480 47.505 207.405 ;
        RECT 47.790 207.245 47.960 207.825 ;
        RECT 48.690 207.405 49.150 207.635 ;
        RECT 48.380 207.260 48.550 207.265 ;
        RECT 47.760 206.595 47.990 207.245 ;
        RECT 48.335 207.230 48.595 207.260 ;
        RECT 48.305 206.970 48.625 207.230 ;
        RECT 48.335 206.940 48.595 206.970 ;
        RECT 48.350 206.595 48.580 206.940 ;
        RECT 47.790 206.575 47.960 206.595 ;
        RECT 47.290 206.435 47.550 206.480 ;
        RECT 47.190 206.205 47.650 206.435 ;
        RECT 47.290 206.160 47.550 206.205 ;
        RECT 47.190 204.270 47.650 204.500 ;
        RECT 46.260 203.065 46.490 204.065 ;
        RECT 46.850 203.360 47.080 204.065 ;
        RECT 46.805 203.100 47.125 203.360 ;
        RECT 46.850 203.065 47.080 203.100 ;
        RECT 45.690 202.830 46.150 202.860 ;
        RECT 45.210 202.660 46.150 202.830 ;
        RECT 45.210 202.615 45.530 202.660 ;
        RECT 45.690 202.630 46.150 202.660 ;
        RECT 46.290 202.470 46.460 203.065 ;
        RECT 46.880 203.045 47.050 203.065 ;
        RECT 46.710 202.830 47.030 202.875 ;
        RECT 47.335 202.860 47.505 204.270 ;
        RECT 47.790 204.065 47.960 204.085 ;
        RECT 48.380 204.065 48.550 206.595 ;
        RECT 48.835 206.480 49.005 207.405 ;
        RECT 49.290 207.245 49.460 207.825 ;
        RECT 50.190 207.405 50.650 207.635 ;
        RECT 49.880 207.260 50.050 207.265 ;
        RECT 49.260 206.595 49.490 207.245 ;
        RECT 49.835 207.230 50.095 207.260 ;
        RECT 49.805 206.970 50.125 207.230 ;
        RECT 49.835 206.940 50.095 206.970 ;
        RECT 49.850 206.595 50.080 206.940 ;
        RECT 49.290 206.575 49.460 206.595 ;
        RECT 48.790 206.435 49.050 206.480 ;
        RECT 48.690 206.205 49.150 206.435 ;
        RECT 48.790 206.160 49.050 206.205 ;
        RECT 48.690 204.270 49.150 204.500 ;
        RECT 47.760 203.065 47.990 204.065 ;
        RECT 48.350 203.360 48.580 204.065 ;
        RECT 48.305 203.100 48.625 203.360 ;
        RECT 48.350 203.065 48.580 203.100 ;
        RECT 47.190 202.830 47.650 202.860 ;
        RECT 46.710 202.660 47.650 202.830 ;
        RECT 46.710 202.615 47.030 202.660 ;
        RECT 47.190 202.630 47.650 202.660 ;
        RECT 47.790 202.470 47.960 203.065 ;
        RECT 48.380 203.045 48.550 203.065 ;
        RECT 48.210 202.830 48.530 202.875 ;
        RECT 48.835 202.860 49.005 204.270 ;
        RECT 49.290 204.065 49.460 204.085 ;
        RECT 49.880 204.065 50.050 206.595 ;
        RECT 50.335 206.480 50.505 207.405 ;
        RECT 50.790 207.245 50.960 207.825 ;
        RECT 51.390 207.810 51.680 207.840 ;
        RECT 64.610 208.130 64.900 208.160 ;
        RECT 66.250 208.130 66.510 208.145 ;
        RECT 67.750 208.130 68.010 208.145 ;
        RECT 69.250 208.130 69.510 208.145 ;
        RECT 70.750 208.130 71.010 208.145 ;
        RECT 72.250 208.130 72.510 208.145 ;
        RECT 73.750 208.130 74.010 208.145 ;
        RECT 75.250 208.130 75.510 208.145 ;
        RECT 76.750 208.130 77.010 208.145 ;
        RECT 77.390 208.130 77.680 208.160 ;
        RECT 64.610 207.840 77.680 208.130 ;
        RECT 64.610 207.810 64.900 207.840 ;
        RECT 66.250 207.825 66.510 207.840 ;
        RECT 67.750 207.825 68.010 207.840 ;
        RECT 69.250 207.825 69.510 207.840 ;
        RECT 70.750 207.825 71.010 207.840 ;
        RECT 72.250 207.825 72.510 207.840 ;
        RECT 73.750 207.825 74.010 207.840 ;
        RECT 75.250 207.825 75.510 207.840 ;
        RECT 76.750 207.825 77.010 207.840 ;
        RECT 65.690 207.405 66.150 207.635 ;
        RECT 65.380 207.260 65.550 207.265 ;
        RECT 50.760 206.595 50.990 207.245 ;
        RECT 65.335 207.230 65.595 207.260 ;
        RECT 65.305 206.970 65.625 207.230 ;
        RECT 65.335 206.940 65.595 206.970 ;
        RECT 65.350 206.595 65.580 206.940 ;
        RECT 50.790 206.575 50.960 206.595 ;
        RECT 50.290 206.435 50.550 206.480 ;
        RECT 50.190 206.205 50.650 206.435 ;
        RECT 50.290 206.160 50.550 206.205 ;
        RECT 50.190 204.270 50.650 204.500 ;
        RECT 49.260 203.065 49.490 204.065 ;
        RECT 49.850 203.360 50.080 204.065 ;
        RECT 49.805 203.100 50.125 203.360 ;
        RECT 49.850 203.065 50.080 203.100 ;
        RECT 48.690 202.830 49.150 202.860 ;
        RECT 48.210 202.660 49.150 202.830 ;
        RECT 48.210 202.615 48.530 202.660 ;
        RECT 48.690 202.630 49.150 202.660 ;
        RECT 49.290 202.470 49.460 203.065 ;
        RECT 49.880 203.045 50.050 203.065 ;
        RECT 49.710 202.830 50.030 202.875 ;
        RECT 50.335 202.860 50.505 204.270 ;
        RECT 50.790 204.065 50.960 204.085 ;
        RECT 65.380 204.065 65.550 206.595 ;
        RECT 65.835 206.480 66.005 207.405 ;
        RECT 66.290 207.245 66.460 207.825 ;
        RECT 67.190 207.405 67.650 207.635 ;
        RECT 66.880 207.260 67.050 207.265 ;
        RECT 66.260 206.595 66.490 207.245 ;
        RECT 66.835 207.230 67.095 207.260 ;
        RECT 66.805 206.970 67.125 207.230 ;
        RECT 66.835 206.940 67.095 206.970 ;
        RECT 66.850 206.595 67.080 206.940 ;
        RECT 66.290 206.575 66.460 206.595 ;
        RECT 65.790 206.435 66.050 206.480 ;
        RECT 65.690 206.205 66.150 206.435 ;
        RECT 65.790 206.160 66.050 206.205 ;
        RECT 65.690 204.270 66.150 204.500 ;
        RECT 50.760 203.065 50.990 204.065 ;
        RECT 65.350 203.360 65.580 204.065 ;
        RECT 65.305 203.100 65.625 203.360 ;
        RECT 65.350 203.065 65.580 203.100 ;
        RECT 50.190 202.830 50.650 202.860 ;
        RECT 49.710 202.660 50.650 202.830 ;
        RECT 49.710 202.615 50.030 202.660 ;
        RECT 50.190 202.630 50.650 202.660 ;
        RECT 50.790 202.470 50.960 203.065 ;
        RECT 65.380 203.045 65.550 203.065 ;
        RECT 65.210 202.830 65.530 202.875 ;
        RECT 65.835 202.860 66.005 204.270 ;
        RECT 66.290 204.065 66.460 204.085 ;
        RECT 66.880 204.065 67.050 206.595 ;
        RECT 67.335 206.480 67.505 207.405 ;
        RECT 67.790 207.245 67.960 207.825 ;
        RECT 68.690 207.405 69.150 207.635 ;
        RECT 68.380 207.260 68.550 207.265 ;
        RECT 67.760 206.595 67.990 207.245 ;
        RECT 68.335 207.230 68.595 207.260 ;
        RECT 68.305 206.970 68.625 207.230 ;
        RECT 68.335 206.940 68.595 206.970 ;
        RECT 68.350 206.595 68.580 206.940 ;
        RECT 67.790 206.575 67.960 206.595 ;
        RECT 67.290 206.435 67.550 206.480 ;
        RECT 67.190 206.205 67.650 206.435 ;
        RECT 67.290 206.160 67.550 206.205 ;
        RECT 67.190 204.270 67.650 204.500 ;
        RECT 66.260 203.065 66.490 204.065 ;
        RECT 66.850 203.360 67.080 204.065 ;
        RECT 66.805 203.100 67.125 203.360 ;
        RECT 66.850 203.065 67.080 203.100 ;
        RECT 65.690 202.830 66.150 202.860 ;
        RECT 65.210 202.660 66.150 202.830 ;
        RECT 65.210 202.615 65.530 202.660 ;
        RECT 65.690 202.630 66.150 202.660 ;
        RECT 51.260 202.470 51.610 202.530 ;
        RECT 13.380 202.290 13.550 202.310 ;
        RECT 13.350 201.640 13.580 202.290 ;
        RECT 13.835 202.050 14.005 202.450 ;
        RECT 14.290 202.290 14.460 202.310 ;
        RECT 14.880 202.290 15.050 202.310 ;
        RECT 14.260 202.050 14.490 202.290 ;
        RECT 13.835 201.880 14.490 202.050 ;
        RECT 13.380 201.060 13.550 201.640 ;
        RECT 13.835 201.480 14.005 201.880 ;
        RECT 14.260 201.640 14.490 201.880 ;
        RECT 14.850 201.640 15.080 202.290 ;
        RECT 15.335 202.050 15.505 202.450 ;
        RECT 15.790 202.290 15.960 202.310 ;
        RECT 16.380 202.290 16.550 202.310 ;
        RECT 15.760 202.050 15.990 202.290 ;
        RECT 15.335 201.880 15.990 202.050 ;
        RECT 14.290 201.620 14.460 201.640 ;
        RECT 13.690 201.250 14.150 201.480 ;
        RECT 14.880 201.060 15.050 201.640 ;
        RECT 15.335 201.480 15.505 201.880 ;
        RECT 15.760 201.640 15.990 201.880 ;
        RECT 16.350 201.640 16.580 202.290 ;
        RECT 16.835 202.050 17.005 202.450 ;
        RECT 17.290 202.290 17.460 202.310 ;
        RECT 17.880 202.290 18.050 202.310 ;
        RECT 17.260 202.050 17.490 202.290 ;
        RECT 16.835 201.880 17.490 202.050 ;
        RECT 15.790 201.620 15.960 201.640 ;
        RECT 15.190 201.250 15.650 201.480 ;
        RECT 16.380 201.060 16.550 201.640 ;
        RECT 16.835 201.480 17.005 201.880 ;
        RECT 17.260 201.640 17.490 201.880 ;
        RECT 17.850 201.640 18.080 202.290 ;
        RECT 18.335 202.050 18.505 202.450 ;
        RECT 18.790 202.290 18.960 202.310 ;
        RECT 19.380 202.290 19.550 202.310 ;
        RECT 18.760 202.050 18.990 202.290 ;
        RECT 18.335 201.880 18.990 202.050 ;
        RECT 17.290 201.620 17.460 201.640 ;
        RECT 16.690 201.250 17.150 201.480 ;
        RECT 17.880 201.060 18.050 201.640 ;
        RECT 18.335 201.480 18.505 201.880 ;
        RECT 18.760 201.640 18.990 201.880 ;
        RECT 19.350 201.640 19.580 202.290 ;
        RECT 19.835 202.050 20.005 202.450 ;
        RECT 20.290 202.290 20.460 202.310 ;
        RECT 20.880 202.290 21.050 202.310 ;
        RECT 20.260 202.050 20.490 202.290 ;
        RECT 19.835 201.880 20.490 202.050 ;
        RECT 18.790 201.620 18.960 201.640 ;
        RECT 18.190 201.250 18.650 201.480 ;
        RECT 19.380 201.060 19.550 201.640 ;
        RECT 19.835 201.480 20.005 201.880 ;
        RECT 20.260 201.640 20.490 201.880 ;
        RECT 20.850 201.640 21.080 202.290 ;
        RECT 21.335 202.050 21.505 202.450 ;
        RECT 21.790 202.290 21.960 202.310 ;
        RECT 22.380 202.290 22.550 202.310 ;
        RECT 21.760 202.050 21.990 202.290 ;
        RECT 21.335 201.880 21.990 202.050 ;
        RECT 20.290 201.620 20.460 201.640 ;
        RECT 19.690 201.250 20.150 201.480 ;
        RECT 20.880 201.060 21.050 201.640 ;
        RECT 21.335 201.480 21.505 201.880 ;
        RECT 21.760 201.640 21.990 201.880 ;
        RECT 22.350 201.640 22.580 202.290 ;
        RECT 22.835 202.050 23.005 202.450 ;
        RECT 23.290 202.290 23.460 202.310 ;
        RECT 23.880 202.290 24.050 202.310 ;
        RECT 23.260 202.050 23.490 202.290 ;
        RECT 22.835 201.880 23.490 202.050 ;
        RECT 21.790 201.620 21.960 201.640 ;
        RECT 21.190 201.250 21.650 201.480 ;
        RECT 22.380 201.060 22.550 201.640 ;
        RECT 22.835 201.480 23.005 201.880 ;
        RECT 23.260 201.640 23.490 201.880 ;
        RECT 23.850 201.640 24.080 202.290 ;
        RECT 24.335 202.050 24.505 202.450 ;
        RECT 24.790 202.290 24.960 202.310 ;
        RECT 24.760 202.050 24.990 202.290 ;
        RECT 38.725 202.180 51.610 202.470 ;
        RECT 38.725 202.120 39.075 202.180 ;
        RECT 51.260 202.120 51.610 202.180 ;
        RECT 64.725 202.470 65.075 202.530 ;
        RECT 66.290 202.470 66.460 203.065 ;
        RECT 66.880 203.045 67.050 203.065 ;
        RECT 66.710 202.830 67.030 202.875 ;
        RECT 67.335 202.860 67.505 204.270 ;
        RECT 67.790 204.065 67.960 204.085 ;
        RECT 68.380 204.065 68.550 206.595 ;
        RECT 68.835 206.480 69.005 207.405 ;
        RECT 69.290 207.245 69.460 207.825 ;
        RECT 70.190 207.405 70.650 207.635 ;
        RECT 69.880 207.260 70.050 207.265 ;
        RECT 69.260 206.595 69.490 207.245 ;
        RECT 69.835 207.230 70.095 207.260 ;
        RECT 69.805 206.970 70.125 207.230 ;
        RECT 69.835 206.940 70.095 206.970 ;
        RECT 69.850 206.595 70.080 206.940 ;
        RECT 69.290 206.575 69.460 206.595 ;
        RECT 68.790 206.435 69.050 206.480 ;
        RECT 68.690 206.205 69.150 206.435 ;
        RECT 68.790 206.160 69.050 206.205 ;
        RECT 68.690 204.270 69.150 204.500 ;
        RECT 67.760 203.065 67.990 204.065 ;
        RECT 68.350 203.360 68.580 204.065 ;
        RECT 68.305 203.100 68.625 203.360 ;
        RECT 68.350 203.065 68.580 203.100 ;
        RECT 67.190 202.830 67.650 202.860 ;
        RECT 66.710 202.660 67.650 202.830 ;
        RECT 66.710 202.615 67.030 202.660 ;
        RECT 67.190 202.630 67.650 202.660 ;
        RECT 67.790 202.470 67.960 203.065 ;
        RECT 68.380 203.045 68.550 203.065 ;
        RECT 68.210 202.830 68.530 202.875 ;
        RECT 68.835 202.860 69.005 204.270 ;
        RECT 69.290 204.065 69.460 204.085 ;
        RECT 69.880 204.065 70.050 206.595 ;
        RECT 70.335 206.480 70.505 207.405 ;
        RECT 70.790 207.245 70.960 207.825 ;
        RECT 71.690 207.405 72.150 207.635 ;
        RECT 71.380 207.260 71.550 207.265 ;
        RECT 70.760 206.595 70.990 207.245 ;
        RECT 71.335 207.230 71.595 207.260 ;
        RECT 71.305 206.970 71.625 207.230 ;
        RECT 71.335 206.940 71.595 206.970 ;
        RECT 71.350 206.595 71.580 206.940 ;
        RECT 70.790 206.575 70.960 206.595 ;
        RECT 70.290 206.435 70.550 206.480 ;
        RECT 70.190 206.205 70.650 206.435 ;
        RECT 70.290 206.160 70.550 206.205 ;
        RECT 70.190 204.270 70.650 204.500 ;
        RECT 69.260 203.065 69.490 204.065 ;
        RECT 69.850 203.360 70.080 204.065 ;
        RECT 69.805 203.100 70.125 203.360 ;
        RECT 69.850 203.065 70.080 203.100 ;
        RECT 68.690 202.830 69.150 202.860 ;
        RECT 68.210 202.660 69.150 202.830 ;
        RECT 68.210 202.615 68.530 202.660 ;
        RECT 68.690 202.630 69.150 202.660 ;
        RECT 69.290 202.470 69.460 203.065 ;
        RECT 69.880 203.045 70.050 203.065 ;
        RECT 69.710 202.830 70.030 202.875 ;
        RECT 70.335 202.860 70.505 204.270 ;
        RECT 70.790 204.065 70.960 204.085 ;
        RECT 71.380 204.065 71.550 206.595 ;
        RECT 71.835 206.480 72.005 207.405 ;
        RECT 72.290 207.245 72.460 207.825 ;
        RECT 73.190 207.405 73.650 207.635 ;
        RECT 72.880 207.260 73.050 207.265 ;
        RECT 72.260 206.595 72.490 207.245 ;
        RECT 72.835 207.230 73.095 207.260 ;
        RECT 72.805 206.970 73.125 207.230 ;
        RECT 72.835 206.940 73.095 206.970 ;
        RECT 72.850 206.595 73.080 206.940 ;
        RECT 72.290 206.575 72.460 206.595 ;
        RECT 71.790 206.435 72.050 206.480 ;
        RECT 71.690 206.205 72.150 206.435 ;
        RECT 71.790 206.160 72.050 206.205 ;
        RECT 71.690 204.270 72.150 204.500 ;
        RECT 70.760 203.065 70.990 204.065 ;
        RECT 71.350 203.360 71.580 204.065 ;
        RECT 71.305 203.100 71.625 203.360 ;
        RECT 71.350 203.065 71.580 203.100 ;
        RECT 70.190 202.830 70.650 202.860 ;
        RECT 69.710 202.660 70.650 202.830 ;
        RECT 69.710 202.615 70.030 202.660 ;
        RECT 70.190 202.630 70.650 202.660 ;
        RECT 70.790 202.470 70.960 203.065 ;
        RECT 71.380 203.045 71.550 203.065 ;
        RECT 71.210 202.830 71.530 202.875 ;
        RECT 71.835 202.860 72.005 204.270 ;
        RECT 72.290 204.065 72.460 204.085 ;
        RECT 72.880 204.065 73.050 206.595 ;
        RECT 73.335 206.480 73.505 207.405 ;
        RECT 73.790 207.245 73.960 207.825 ;
        RECT 74.690 207.405 75.150 207.635 ;
        RECT 74.380 207.260 74.550 207.265 ;
        RECT 73.760 206.595 73.990 207.245 ;
        RECT 74.335 207.230 74.595 207.260 ;
        RECT 74.305 206.970 74.625 207.230 ;
        RECT 74.335 206.940 74.595 206.970 ;
        RECT 74.350 206.595 74.580 206.940 ;
        RECT 73.790 206.575 73.960 206.595 ;
        RECT 73.290 206.435 73.550 206.480 ;
        RECT 73.190 206.205 73.650 206.435 ;
        RECT 73.290 206.160 73.550 206.205 ;
        RECT 73.190 204.270 73.650 204.500 ;
        RECT 72.260 203.065 72.490 204.065 ;
        RECT 72.850 203.360 73.080 204.065 ;
        RECT 72.805 203.100 73.125 203.360 ;
        RECT 72.850 203.065 73.080 203.100 ;
        RECT 71.690 202.830 72.150 202.860 ;
        RECT 71.210 202.660 72.150 202.830 ;
        RECT 71.210 202.615 71.530 202.660 ;
        RECT 71.690 202.630 72.150 202.660 ;
        RECT 72.290 202.470 72.460 203.065 ;
        RECT 72.880 203.045 73.050 203.065 ;
        RECT 72.710 202.830 73.030 202.875 ;
        RECT 73.335 202.860 73.505 204.270 ;
        RECT 73.790 204.065 73.960 204.085 ;
        RECT 74.380 204.065 74.550 206.595 ;
        RECT 74.835 206.480 75.005 207.405 ;
        RECT 75.290 207.245 75.460 207.825 ;
        RECT 76.190 207.405 76.650 207.635 ;
        RECT 75.880 207.260 76.050 207.265 ;
        RECT 75.260 206.595 75.490 207.245 ;
        RECT 75.835 207.230 76.095 207.260 ;
        RECT 75.805 206.970 76.125 207.230 ;
        RECT 75.835 206.940 76.095 206.970 ;
        RECT 75.850 206.595 76.080 206.940 ;
        RECT 75.290 206.575 75.460 206.595 ;
        RECT 74.790 206.435 75.050 206.480 ;
        RECT 74.690 206.205 75.150 206.435 ;
        RECT 74.790 206.160 75.050 206.205 ;
        RECT 74.690 204.270 75.150 204.500 ;
        RECT 73.760 203.065 73.990 204.065 ;
        RECT 74.350 203.360 74.580 204.065 ;
        RECT 74.305 203.100 74.625 203.360 ;
        RECT 74.350 203.065 74.580 203.100 ;
        RECT 73.190 202.830 73.650 202.860 ;
        RECT 72.710 202.660 73.650 202.830 ;
        RECT 72.710 202.615 73.030 202.660 ;
        RECT 73.190 202.630 73.650 202.660 ;
        RECT 73.790 202.470 73.960 203.065 ;
        RECT 74.380 203.045 74.550 203.065 ;
        RECT 74.210 202.830 74.530 202.875 ;
        RECT 74.835 202.860 75.005 204.270 ;
        RECT 75.290 204.065 75.460 204.085 ;
        RECT 75.880 204.065 76.050 206.595 ;
        RECT 76.335 206.480 76.505 207.405 ;
        RECT 76.790 207.245 76.960 207.825 ;
        RECT 77.390 207.810 77.680 207.840 ;
        RECT 76.760 206.595 76.990 207.245 ;
        RECT 106.760 206.625 107.050 206.655 ;
        RECT 107.265 206.625 107.525 206.640 ;
        RECT 108.765 206.625 109.025 206.640 ;
        RECT 110.265 206.625 110.525 206.640 ;
        RECT 111.765 206.625 112.025 206.640 ;
        RECT 113.265 206.625 113.525 206.640 ;
        RECT 114.765 206.625 115.025 206.640 ;
        RECT 116.265 206.625 116.525 206.640 ;
        RECT 117.765 206.625 118.025 206.640 ;
        RECT 119.290 206.625 119.580 206.655 ;
        RECT 76.790 206.575 76.960 206.595 ;
        RECT 76.290 206.435 76.550 206.480 ;
        RECT 76.190 206.205 76.650 206.435 ;
        RECT 106.760 206.335 119.580 206.625 ;
        RECT 106.760 206.305 107.050 206.335 ;
        RECT 107.265 206.320 107.550 206.335 ;
        RECT 108.765 206.320 109.050 206.335 ;
        RECT 110.265 206.320 110.550 206.335 ;
        RECT 111.765 206.320 112.050 206.335 ;
        RECT 113.265 206.320 113.550 206.335 ;
        RECT 114.765 206.320 115.050 206.335 ;
        RECT 116.265 206.320 116.550 206.335 ;
        RECT 117.765 206.320 118.050 206.335 ;
        RECT 76.290 206.160 76.550 206.205 ;
        RECT 107.380 205.740 107.550 206.320 ;
        RECT 107.690 205.945 108.150 206.175 ;
        RECT 107.760 205.805 108.080 205.945 ;
        RECT 107.350 204.740 107.580 205.740 ;
        RECT 107.380 204.720 107.550 204.740 ;
        RECT 107.835 204.535 108.005 205.805 ;
        RECT 108.290 205.740 108.460 205.760 ;
        RECT 108.880 205.740 109.050 206.320 ;
        RECT 109.190 205.945 109.650 206.175 ;
        RECT 109.260 205.805 109.580 205.945 ;
        RECT 108.260 204.740 108.490 205.740 ;
        RECT 108.850 204.740 109.080 205.740 ;
        RECT 76.190 204.270 76.650 204.500 ;
        RECT 107.690 204.305 108.150 204.535 ;
        RECT 75.260 203.065 75.490 204.065 ;
        RECT 75.850 203.360 76.080 204.065 ;
        RECT 75.805 203.100 76.125 203.360 ;
        RECT 75.850 203.065 76.080 203.100 ;
        RECT 74.690 202.830 75.150 202.860 ;
        RECT 74.210 202.660 75.150 202.830 ;
        RECT 74.210 202.615 74.530 202.660 ;
        RECT 74.690 202.630 75.150 202.660 ;
        RECT 75.290 202.470 75.460 203.065 ;
        RECT 75.880 203.045 76.050 203.065 ;
        RECT 75.710 202.830 76.030 202.875 ;
        RECT 76.335 202.860 76.505 204.270 ;
        RECT 76.790 204.065 76.960 204.085 ;
        RECT 76.760 203.065 76.990 204.065 ;
        RECT 76.190 202.830 76.650 202.860 ;
        RECT 75.710 202.660 76.650 202.830 ;
        RECT 75.710 202.615 76.030 202.660 ;
        RECT 76.190 202.630 76.650 202.660 ;
        RECT 76.790 202.470 76.960 203.065 ;
        RECT 107.835 202.600 108.005 204.305 ;
        RECT 77.260 202.470 77.610 202.530 ;
        RECT 64.725 202.180 77.610 202.470 ;
        RECT 107.690 202.370 108.150 202.600 ;
        RECT 107.380 202.210 107.550 202.230 ;
        RECT 64.725 202.120 65.075 202.180 ;
        RECT 77.260 202.120 77.610 202.180 ;
        RECT 24.335 201.880 24.990 202.050 ;
        RECT 23.290 201.620 23.460 201.640 ;
        RECT 22.690 201.250 23.150 201.480 ;
        RECT 23.880 201.060 24.050 201.640 ;
        RECT 24.335 201.480 24.505 201.880 ;
        RECT 24.760 201.640 24.990 201.880 ;
        RECT 24.790 201.620 24.960 201.640 ;
        RECT 107.350 201.560 107.580 202.210 ;
        RECT 24.190 201.250 24.650 201.480 ;
        RECT 38.580 201.420 38.930 201.480 ;
        RECT 51.360 201.420 51.710 201.480 ;
        RECT 38.580 201.130 51.710 201.420 ;
        RECT 38.580 201.070 38.930 201.130 ;
        RECT 13.335 201.045 13.595 201.060 ;
        RECT 14.835 201.045 15.095 201.060 ;
        RECT 16.335 201.045 16.595 201.060 ;
        RECT 17.835 201.045 18.095 201.060 ;
        RECT 19.335 201.045 19.595 201.060 ;
        RECT 20.835 201.045 21.095 201.060 ;
        RECT 22.335 201.045 22.595 201.060 ;
        RECT 23.835 201.045 24.095 201.060 ;
        RECT 13.170 200.755 25.170 201.045 ;
        RECT 13.335 200.740 13.595 200.755 ;
        RECT 14.835 200.740 15.095 200.755 ;
        RECT 16.335 200.740 16.595 200.755 ;
        RECT 17.835 200.740 18.095 200.755 ;
        RECT 19.335 200.740 19.595 200.755 ;
        RECT 20.835 200.740 21.095 200.755 ;
        RECT 22.335 200.740 22.595 200.755 ;
        RECT 23.835 200.740 24.095 200.755 ;
        RECT 39.690 200.695 40.150 200.925 ;
        RECT 39.380 200.550 39.550 200.555 ;
        RECT 39.335 200.230 39.595 200.550 ;
        RECT 39.350 199.885 39.580 200.230 ;
        RECT 39.380 197.355 39.550 199.885 ;
        RECT 39.835 199.725 40.005 200.695 ;
        RECT 40.290 200.535 40.460 201.130 ;
        RECT 41.190 200.695 41.650 200.925 ;
        RECT 40.880 200.550 41.050 200.555 ;
        RECT 40.260 199.885 40.490 200.535 ;
        RECT 40.835 200.230 41.095 200.550 ;
        RECT 40.850 199.885 41.080 200.230 ;
        RECT 40.290 199.865 40.460 199.885 ;
        RECT 39.690 199.695 40.150 199.725 ;
        RECT 39.690 199.525 40.460 199.695 ;
        RECT 39.690 199.495 40.150 199.525 ;
        RECT 39.760 199.075 40.080 199.335 ;
        RECT 39.835 197.835 40.005 199.075 ;
        RECT 40.290 198.445 40.460 199.525 ;
        RECT 40.245 198.125 40.505 198.445 ;
        RECT 39.790 197.790 40.050 197.835 ;
        RECT 39.690 197.560 40.150 197.790 ;
        RECT 39.790 197.515 40.050 197.560 ;
        RECT 39.350 196.355 39.580 197.355 ;
        RECT 39.380 196.335 39.550 196.355 ;
        RECT 39.835 196.150 40.005 197.515 ;
        RECT 40.290 197.355 40.460 197.375 ;
        RECT 40.880 197.355 41.050 199.885 ;
        RECT 41.335 199.725 41.505 200.695 ;
        RECT 41.790 200.535 41.960 201.130 ;
        RECT 42.690 200.695 43.150 200.925 ;
        RECT 42.380 200.550 42.550 200.555 ;
        RECT 41.760 199.885 41.990 200.535 ;
        RECT 42.335 200.230 42.595 200.550 ;
        RECT 42.350 199.885 42.580 200.230 ;
        RECT 41.790 199.865 41.960 199.885 ;
        RECT 41.190 199.695 41.650 199.725 ;
        RECT 41.190 199.525 41.960 199.695 ;
        RECT 41.190 199.495 41.650 199.525 ;
        RECT 41.260 199.075 41.580 199.335 ;
        RECT 41.335 197.835 41.505 199.075 ;
        RECT 41.790 198.445 41.960 199.525 ;
        RECT 41.745 198.125 42.005 198.445 ;
        RECT 41.290 197.790 41.550 197.835 ;
        RECT 41.190 197.560 41.650 197.790 ;
        RECT 41.290 197.515 41.550 197.560 ;
        RECT 40.260 196.355 40.490 197.355 ;
        RECT 40.850 196.355 41.080 197.355 ;
        RECT 39.690 195.920 40.150 196.150 ;
        RECT 38.760 195.760 39.050 195.790 ;
        RECT 40.290 195.775 40.460 196.355 ;
        RECT 40.880 196.335 41.050 196.355 ;
        RECT 41.335 196.150 41.505 197.515 ;
        RECT 41.790 197.355 41.960 197.375 ;
        RECT 42.380 197.355 42.550 199.885 ;
        RECT 42.835 199.725 43.005 200.695 ;
        RECT 43.290 200.535 43.460 201.130 ;
        RECT 44.190 200.695 44.650 200.925 ;
        RECT 43.880 200.550 44.050 200.555 ;
        RECT 43.260 199.885 43.490 200.535 ;
        RECT 43.835 200.230 44.095 200.550 ;
        RECT 43.850 199.885 44.080 200.230 ;
        RECT 43.290 199.865 43.460 199.885 ;
        RECT 42.690 199.695 43.150 199.725 ;
        RECT 42.690 199.525 43.460 199.695 ;
        RECT 42.690 199.495 43.150 199.525 ;
        RECT 42.760 199.075 43.080 199.335 ;
        RECT 42.835 197.835 43.005 199.075 ;
        RECT 43.290 198.445 43.460 199.525 ;
        RECT 43.245 198.125 43.505 198.445 ;
        RECT 42.790 197.790 43.050 197.835 ;
        RECT 42.690 197.560 43.150 197.790 ;
        RECT 42.790 197.515 43.050 197.560 ;
        RECT 41.760 196.355 41.990 197.355 ;
        RECT 42.350 196.355 42.580 197.355 ;
        RECT 41.190 195.920 41.650 196.150 ;
        RECT 41.790 195.775 41.960 196.355 ;
        RECT 42.380 196.335 42.550 196.355 ;
        RECT 42.835 196.150 43.005 197.515 ;
        RECT 43.290 197.355 43.460 197.375 ;
        RECT 43.880 197.355 44.050 199.885 ;
        RECT 44.335 199.725 44.505 200.695 ;
        RECT 44.790 200.535 44.960 201.130 ;
        RECT 45.690 200.695 46.150 200.925 ;
        RECT 45.380 200.550 45.550 200.555 ;
        RECT 44.760 199.885 44.990 200.535 ;
        RECT 45.335 200.230 45.595 200.550 ;
        RECT 45.350 199.885 45.580 200.230 ;
        RECT 44.790 199.865 44.960 199.885 ;
        RECT 44.190 199.695 44.650 199.725 ;
        RECT 44.190 199.525 44.960 199.695 ;
        RECT 44.190 199.495 44.650 199.525 ;
        RECT 44.260 199.075 44.580 199.335 ;
        RECT 44.335 197.835 44.505 199.075 ;
        RECT 44.790 198.445 44.960 199.525 ;
        RECT 44.745 198.125 45.005 198.445 ;
        RECT 44.290 197.790 44.550 197.835 ;
        RECT 44.190 197.560 44.650 197.790 ;
        RECT 44.290 197.515 44.550 197.560 ;
        RECT 43.260 196.355 43.490 197.355 ;
        RECT 43.850 196.355 44.080 197.355 ;
        RECT 42.690 195.920 43.150 196.150 ;
        RECT 43.290 195.775 43.460 196.355 ;
        RECT 43.880 196.335 44.050 196.355 ;
        RECT 44.335 196.150 44.505 197.515 ;
        RECT 44.790 197.355 44.960 197.375 ;
        RECT 45.380 197.355 45.550 199.885 ;
        RECT 45.835 199.725 46.005 200.695 ;
        RECT 46.290 200.535 46.460 201.130 ;
        RECT 47.190 200.695 47.650 200.925 ;
        RECT 46.880 200.550 47.050 200.555 ;
        RECT 46.260 199.885 46.490 200.535 ;
        RECT 46.835 200.230 47.095 200.550 ;
        RECT 46.850 199.885 47.080 200.230 ;
        RECT 46.290 199.865 46.460 199.885 ;
        RECT 45.690 199.695 46.150 199.725 ;
        RECT 45.690 199.525 46.460 199.695 ;
        RECT 45.690 199.495 46.150 199.525 ;
        RECT 45.760 199.075 46.080 199.335 ;
        RECT 45.835 197.835 46.005 199.075 ;
        RECT 46.290 198.445 46.460 199.525 ;
        RECT 46.245 198.125 46.505 198.445 ;
        RECT 45.790 197.790 46.050 197.835 ;
        RECT 45.690 197.560 46.150 197.790 ;
        RECT 45.790 197.515 46.050 197.560 ;
        RECT 44.760 196.355 44.990 197.355 ;
        RECT 45.350 196.355 45.580 197.355 ;
        RECT 44.190 195.920 44.650 196.150 ;
        RECT 44.790 195.775 44.960 196.355 ;
        RECT 45.380 196.335 45.550 196.355 ;
        RECT 45.835 196.150 46.005 197.515 ;
        RECT 46.290 197.355 46.460 197.375 ;
        RECT 46.880 197.355 47.050 199.885 ;
        RECT 47.335 199.725 47.505 200.695 ;
        RECT 47.790 200.535 47.960 201.130 ;
        RECT 48.690 200.695 49.150 200.925 ;
        RECT 48.380 200.550 48.550 200.555 ;
        RECT 47.760 199.885 47.990 200.535 ;
        RECT 48.335 200.230 48.595 200.550 ;
        RECT 48.350 199.885 48.580 200.230 ;
        RECT 47.790 199.865 47.960 199.885 ;
        RECT 47.190 199.695 47.650 199.725 ;
        RECT 47.190 199.525 47.960 199.695 ;
        RECT 47.190 199.495 47.650 199.525 ;
        RECT 47.260 199.075 47.580 199.335 ;
        RECT 47.335 197.835 47.505 199.075 ;
        RECT 47.790 198.445 47.960 199.525 ;
        RECT 47.745 198.125 48.005 198.445 ;
        RECT 47.290 197.790 47.550 197.835 ;
        RECT 47.190 197.560 47.650 197.790 ;
        RECT 47.290 197.515 47.550 197.560 ;
        RECT 46.260 196.355 46.490 197.355 ;
        RECT 46.850 196.355 47.080 197.355 ;
        RECT 45.690 195.920 46.150 196.150 ;
        RECT 46.290 195.775 46.460 196.355 ;
        RECT 46.880 196.335 47.050 196.355 ;
        RECT 47.335 196.150 47.505 197.515 ;
        RECT 47.790 197.355 47.960 197.375 ;
        RECT 48.380 197.355 48.550 199.885 ;
        RECT 48.835 199.725 49.005 200.695 ;
        RECT 49.290 200.535 49.460 201.130 ;
        RECT 50.190 200.695 50.650 200.925 ;
        RECT 49.880 200.550 50.050 200.555 ;
        RECT 49.260 199.885 49.490 200.535 ;
        RECT 49.835 200.230 50.095 200.550 ;
        RECT 49.850 199.885 50.080 200.230 ;
        RECT 49.290 199.865 49.460 199.885 ;
        RECT 48.690 199.695 49.150 199.725 ;
        RECT 48.690 199.525 49.460 199.695 ;
        RECT 48.690 199.495 49.150 199.525 ;
        RECT 48.760 199.075 49.080 199.335 ;
        RECT 48.835 197.835 49.005 199.075 ;
        RECT 49.290 198.445 49.460 199.525 ;
        RECT 49.245 198.125 49.505 198.445 ;
        RECT 48.790 197.790 49.050 197.835 ;
        RECT 48.690 197.560 49.150 197.790 ;
        RECT 48.790 197.515 49.050 197.560 ;
        RECT 47.760 196.355 47.990 197.355 ;
        RECT 48.350 196.355 48.580 197.355 ;
        RECT 47.190 195.920 47.650 196.150 ;
        RECT 47.790 195.775 47.960 196.355 ;
        RECT 48.380 196.335 48.550 196.355 ;
        RECT 48.835 196.150 49.005 197.515 ;
        RECT 49.290 197.355 49.460 197.375 ;
        RECT 49.880 197.355 50.050 199.885 ;
        RECT 50.335 199.725 50.505 200.695 ;
        RECT 50.790 200.535 50.960 201.130 ;
        RECT 51.360 201.070 51.710 201.130 ;
        RECT 64.580 201.420 64.930 201.480 ;
        RECT 77.360 201.420 77.710 201.480 ;
        RECT 64.580 201.130 77.710 201.420 ;
        RECT 64.580 201.070 64.930 201.130 ;
        RECT 65.690 200.695 66.150 200.925 ;
        RECT 65.380 200.550 65.550 200.555 ;
        RECT 50.760 199.885 50.990 200.535 ;
        RECT 65.335 200.230 65.595 200.550 ;
        RECT 65.350 199.885 65.580 200.230 ;
        RECT 50.790 199.865 50.960 199.885 ;
        RECT 50.190 199.695 50.650 199.725 ;
        RECT 50.190 199.525 50.960 199.695 ;
        RECT 50.190 199.495 50.650 199.525 ;
        RECT 50.260 199.075 50.580 199.335 ;
        RECT 50.335 197.835 50.505 199.075 ;
        RECT 50.790 198.445 50.960 199.525 ;
        RECT 50.745 198.125 51.005 198.445 ;
        RECT 50.290 197.790 50.550 197.835 ;
        RECT 50.190 197.560 50.650 197.790 ;
        RECT 50.290 197.515 50.550 197.560 ;
        RECT 49.260 196.355 49.490 197.355 ;
        RECT 49.850 196.355 50.080 197.355 ;
        RECT 48.690 195.920 49.150 196.150 ;
        RECT 49.290 195.775 49.460 196.355 ;
        RECT 49.880 196.335 50.050 196.355 ;
        RECT 50.335 196.150 50.505 197.515 ;
        RECT 50.790 197.355 50.960 197.375 ;
        RECT 65.380 197.355 65.550 199.885 ;
        RECT 65.835 199.725 66.005 200.695 ;
        RECT 66.290 200.535 66.460 201.130 ;
        RECT 67.190 200.695 67.650 200.925 ;
        RECT 66.880 200.550 67.050 200.555 ;
        RECT 66.260 199.885 66.490 200.535 ;
        RECT 66.835 200.230 67.095 200.550 ;
        RECT 66.850 199.885 67.080 200.230 ;
        RECT 66.290 199.865 66.460 199.885 ;
        RECT 65.690 199.695 66.150 199.725 ;
        RECT 65.690 199.525 66.460 199.695 ;
        RECT 65.690 199.495 66.150 199.525 ;
        RECT 65.760 199.075 66.080 199.335 ;
        RECT 65.835 197.835 66.005 199.075 ;
        RECT 66.290 198.445 66.460 199.525 ;
        RECT 66.245 198.125 66.505 198.445 ;
        RECT 65.790 197.790 66.050 197.835 ;
        RECT 65.690 197.560 66.150 197.790 ;
        RECT 65.790 197.515 66.050 197.560 ;
        RECT 50.760 196.355 50.990 197.355 ;
        RECT 65.350 196.355 65.580 197.355 ;
        RECT 50.190 195.920 50.650 196.150 ;
        RECT 50.790 195.775 50.960 196.355 ;
        RECT 65.380 196.335 65.550 196.355 ;
        RECT 65.835 196.150 66.005 197.515 ;
        RECT 66.290 197.355 66.460 197.375 ;
        RECT 66.880 197.355 67.050 199.885 ;
        RECT 67.335 199.725 67.505 200.695 ;
        RECT 67.790 200.535 67.960 201.130 ;
        RECT 68.690 200.695 69.150 200.925 ;
        RECT 68.380 200.550 68.550 200.555 ;
        RECT 67.760 199.885 67.990 200.535 ;
        RECT 68.335 200.230 68.595 200.550 ;
        RECT 68.350 199.885 68.580 200.230 ;
        RECT 67.790 199.865 67.960 199.885 ;
        RECT 67.190 199.695 67.650 199.725 ;
        RECT 67.190 199.525 67.960 199.695 ;
        RECT 67.190 199.495 67.650 199.525 ;
        RECT 67.260 199.075 67.580 199.335 ;
        RECT 67.335 197.835 67.505 199.075 ;
        RECT 67.790 198.445 67.960 199.525 ;
        RECT 67.745 198.125 68.005 198.445 ;
        RECT 67.290 197.790 67.550 197.835 ;
        RECT 67.190 197.560 67.650 197.790 ;
        RECT 67.290 197.515 67.550 197.560 ;
        RECT 66.260 196.355 66.490 197.355 ;
        RECT 66.850 196.355 67.080 197.355 ;
        RECT 65.690 195.920 66.150 196.150 ;
        RECT 40.245 195.760 40.505 195.775 ;
        RECT 41.745 195.760 42.005 195.775 ;
        RECT 43.245 195.760 43.505 195.775 ;
        RECT 44.745 195.760 45.005 195.775 ;
        RECT 46.245 195.760 46.505 195.775 ;
        RECT 47.745 195.760 48.005 195.775 ;
        RECT 49.245 195.760 49.505 195.775 ;
        RECT 50.745 195.760 51.005 195.775 ;
        RECT 51.290 195.760 51.580 195.790 ;
        RECT 38.760 195.470 51.580 195.760 ;
        RECT 38.760 195.440 39.050 195.470 ;
        RECT 40.245 195.455 40.505 195.470 ;
        RECT 41.745 195.455 42.005 195.470 ;
        RECT 43.245 195.455 43.505 195.470 ;
        RECT 44.745 195.455 45.005 195.470 ;
        RECT 46.245 195.455 46.505 195.470 ;
        RECT 47.745 195.455 48.005 195.470 ;
        RECT 49.245 195.455 49.505 195.470 ;
        RECT 50.745 195.455 51.005 195.470 ;
        RECT 51.290 195.440 51.580 195.470 ;
        RECT 64.760 195.760 65.050 195.790 ;
        RECT 66.290 195.775 66.460 196.355 ;
        RECT 66.880 196.335 67.050 196.355 ;
        RECT 67.335 196.150 67.505 197.515 ;
        RECT 67.790 197.355 67.960 197.375 ;
        RECT 68.380 197.355 68.550 199.885 ;
        RECT 68.835 199.725 69.005 200.695 ;
        RECT 69.290 200.535 69.460 201.130 ;
        RECT 70.190 200.695 70.650 200.925 ;
        RECT 69.880 200.550 70.050 200.555 ;
        RECT 69.260 199.885 69.490 200.535 ;
        RECT 69.835 200.230 70.095 200.550 ;
        RECT 69.850 199.885 70.080 200.230 ;
        RECT 69.290 199.865 69.460 199.885 ;
        RECT 68.690 199.695 69.150 199.725 ;
        RECT 68.690 199.525 69.460 199.695 ;
        RECT 68.690 199.495 69.150 199.525 ;
        RECT 68.760 199.075 69.080 199.335 ;
        RECT 68.835 197.835 69.005 199.075 ;
        RECT 69.290 198.445 69.460 199.525 ;
        RECT 69.245 198.125 69.505 198.445 ;
        RECT 68.790 197.790 69.050 197.835 ;
        RECT 68.690 197.560 69.150 197.790 ;
        RECT 68.790 197.515 69.050 197.560 ;
        RECT 67.760 196.355 67.990 197.355 ;
        RECT 68.350 196.355 68.580 197.355 ;
        RECT 67.190 195.920 67.650 196.150 ;
        RECT 67.790 195.775 67.960 196.355 ;
        RECT 68.380 196.335 68.550 196.355 ;
        RECT 68.835 196.150 69.005 197.515 ;
        RECT 69.290 197.355 69.460 197.375 ;
        RECT 69.880 197.355 70.050 199.885 ;
        RECT 70.335 199.725 70.505 200.695 ;
        RECT 70.790 200.535 70.960 201.130 ;
        RECT 71.690 200.695 72.150 200.925 ;
        RECT 71.380 200.550 71.550 200.555 ;
        RECT 70.760 199.885 70.990 200.535 ;
        RECT 71.335 200.230 71.595 200.550 ;
        RECT 71.350 199.885 71.580 200.230 ;
        RECT 70.790 199.865 70.960 199.885 ;
        RECT 70.190 199.695 70.650 199.725 ;
        RECT 70.190 199.525 70.960 199.695 ;
        RECT 70.190 199.495 70.650 199.525 ;
        RECT 70.260 199.075 70.580 199.335 ;
        RECT 70.335 197.835 70.505 199.075 ;
        RECT 70.790 198.445 70.960 199.525 ;
        RECT 70.745 198.125 71.005 198.445 ;
        RECT 70.290 197.790 70.550 197.835 ;
        RECT 70.190 197.560 70.650 197.790 ;
        RECT 70.290 197.515 70.550 197.560 ;
        RECT 69.260 196.355 69.490 197.355 ;
        RECT 69.850 196.355 70.080 197.355 ;
        RECT 68.690 195.920 69.150 196.150 ;
        RECT 69.290 195.775 69.460 196.355 ;
        RECT 69.880 196.335 70.050 196.355 ;
        RECT 70.335 196.150 70.505 197.515 ;
        RECT 70.790 197.355 70.960 197.375 ;
        RECT 71.380 197.355 71.550 199.885 ;
        RECT 71.835 199.725 72.005 200.695 ;
        RECT 72.290 200.535 72.460 201.130 ;
        RECT 73.190 200.695 73.650 200.925 ;
        RECT 72.880 200.550 73.050 200.555 ;
        RECT 72.260 199.885 72.490 200.535 ;
        RECT 72.835 200.230 73.095 200.550 ;
        RECT 72.850 199.885 73.080 200.230 ;
        RECT 72.290 199.865 72.460 199.885 ;
        RECT 71.690 199.695 72.150 199.725 ;
        RECT 71.690 199.525 72.460 199.695 ;
        RECT 71.690 199.495 72.150 199.525 ;
        RECT 71.760 199.075 72.080 199.335 ;
        RECT 71.835 197.835 72.005 199.075 ;
        RECT 72.290 198.445 72.460 199.525 ;
        RECT 72.245 198.125 72.505 198.445 ;
        RECT 71.790 197.790 72.050 197.835 ;
        RECT 71.690 197.560 72.150 197.790 ;
        RECT 71.790 197.515 72.050 197.560 ;
        RECT 70.760 196.355 70.990 197.355 ;
        RECT 71.350 196.355 71.580 197.355 ;
        RECT 70.190 195.920 70.650 196.150 ;
        RECT 70.790 195.775 70.960 196.355 ;
        RECT 71.380 196.335 71.550 196.355 ;
        RECT 71.835 196.150 72.005 197.515 ;
        RECT 72.290 197.355 72.460 197.375 ;
        RECT 72.880 197.355 73.050 199.885 ;
        RECT 73.335 199.725 73.505 200.695 ;
        RECT 73.790 200.535 73.960 201.130 ;
        RECT 74.690 200.695 75.150 200.925 ;
        RECT 74.380 200.550 74.550 200.555 ;
        RECT 73.760 199.885 73.990 200.535 ;
        RECT 74.335 200.230 74.595 200.550 ;
        RECT 74.350 199.885 74.580 200.230 ;
        RECT 73.790 199.865 73.960 199.885 ;
        RECT 73.190 199.695 73.650 199.725 ;
        RECT 73.190 199.525 73.960 199.695 ;
        RECT 73.190 199.495 73.650 199.525 ;
        RECT 73.260 199.075 73.580 199.335 ;
        RECT 73.335 197.835 73.505 199.075 ;
        RECT 73.790 198.445 73.960 199.525 ;
        RECT 73.745 198.125 74.005 198.445 ;
        RECT 73.290 197.790 73.550 197.835 ;
        RECT 73.190 197.560 73.650 197.790 ;
        RECT 73.290 197.515 73.550 197.560 ;
        RECT 72.260 196.355 72.490 197.355 ;
        RECT 72.850 196.355 73.080 197.355 ;
        RECT 71.690 195.920 72.150 196.150 ;
        RECT 72.290 195.775 72.460 196.355 ;
        RECT 72.880 196.335 73.050 196.355 ;
        RECT 73.335 196.150 73.505 197.515 ;
        RECT 73.790 197.355 73.960 197.375 ;
        RECT 74.380 197.355 74.550 199.885 ;
        RECT 74.835 199.725 75.005 200.695 ;
        RECT 75.290 200.535 75.460 201.130 ;
        RECT 76.190 200.695 76.650 200.925 ;
        RECT 75.880 200.550 76.050 200.555 ;
        RECT 75.260 199.885 75.490 200.535 ;
        RECT 75.835 200.230 76.095 200.550 ;
        RECT 75.850 199.885 76.080 200.230 ;
        RECT 75.290 199.865 75.460 199.885 ;
        RECT 74.690 199.695 75.150 199.725 ;
        RECT 74.690 199.525 75.460 199.695 ;
        RECT 74.690 199.495 75.150 199.525 ;
        RECT 74.760 199.075 75.080 199.335 ;
        RECT 74.835 197.835 75.005 199.075 ;
        RECT 75.290 198.445 75.460 199.525 ;
        RECT 75.245 198.125 75.505 198.445 ;
        RECT 74.790 197.790 75.050 197.835 ;
        RECT 74.690 197.560 75.150 197.790 ;
        RECT 74.790 197.515 75.050 197.560 ;
        RECT 73.760 196.355 73.990 197.355 ;
        RECT 74.350 196.355 74.580 197.355 ;
        RECT 73.190 195.920 73.650 196.150 ;
        RECT 73.790 195.775 73.960 196.355 ;
        RECT 74.380 196.335 74.550 196.355 ;
        RECT 74.835 196.150 75.005 197.515 ;
        RECT 75.290 197.355 75.460 197.375 ;
        RECT 75.880 197.355 76.050 199.885 ;
        RECT 76.335 199.725 76.505 200.695 ;
        RECT 76.790 200.535 76.960 201.130 ;
        RECT 77.360 201.070 77.710 201.130 ;
        RECT 107.380 200.980 107.550 201.560 ;
        RECT 107.835 201.415 108.005 202.370 ;
        RECT 108.290 202.210 108.460 204.740 ;
        RECT 108.880 204.720 109.050 204.740 ;
        RECT 109.335 204.535 109.505 205.805 ;
        RECT 109.790 205.740 109.960 205.760 ;
        RECT 110.380 205.740 110.550 206.320 ;
        RECT 110.690 205.945 111.150 206.175 ;
        RECT 110.760 205.805 111.080 205.945 ;
        RECT 109.760 204.740 109.990 205.740 ;
        RECT 110.350 204.740 110.580 205.740 ;
        RECT 109.190 204.305 109.650 204.535 ;
        RECT 109.335 202.600 109.505 204.305 ;
        RECT 109.190 202.370 109.650 202.600 ;
        RECT 108.880 202.210 109.050 202.230 ;
        RECT 108.260 201.835 108.490 202.210 ;
        RECT 108.215 201.575 108.535 201.835 ;
        RECT 108.260 201.560 108.490 201.575 ;
        RECT 108.850 201.560 109.080 202.210 ;
        RECT 108.290 201.540 108.460 201.560 ;
        RECT 107.760 201.400 108.080 201.415 ;
        RECT 107.690 201.170 108.150 201.400 ;
        RECT 107.760 201.155 108.080 201.170 ;
        RECT 108.880 200.980 109.050 201.560 ;
        RECT 109.335 201.415 109.505 202.370 ;
        RECT 109.790 202.210 109.960 204.740 ;
        RECT 110.380 204.720 110.550 204.740 ;
        RECT 110.835 204.535 111.005 205.805 ;
        RECT 111.290 205.740 111.460 205.760 ;
        RECT 111.880 205.740 112.050 206.320 ;
        RECT 112.190 205.945 112.650 206.175 ;
        RECT 112.260 205.805 112.580 205.945 ;
        RECT 111.260 204.740 111.490 205.740 ;
        RECT 111.850 204.740 112.080 205.740 ;
        RECT 110.690 204.305 111.150 204.535 ;
        RECT 110.835 202.600 111.005 204.305 ;
        RECT 110.690 202.370 111.150 202.600 ;
        RECT 110.380 202.210 110.550 202.230 ;
        RECT 109.760 201.835 109.990 202.210 ;
        RECT 109.715 201.575 110.035 201.835 ;
        RECT 109.760 201.560 109.990 201.575 ;
        RECT 110.350 201.560 110.580 202.210 ;
        RECT 109.790 201.540 109.960 201.560 ;
        RECT 109.260 201.400 109.580 201.415 ;
        RECT 109.190 201.170 109.650 201.400 ;
        RECT 109.260 201.155 109.580 201.170 ;
        RECT 110.380 200.980 110.550 201.560 ;
        RECT 110.835 201.415 111.005 202.370 ;
        RECT 111.290 202.210 111.460 204.740 ;
        RECT 111.880 204.720 112.050 204.740 ;
        RECT 112.335 204.535 112.505 205.805 ;
        RECT 112.790 205.740 112.960 205.760 ;
        RECT 113.380 205.740 113.550 206.320 ;
        RECT 113.690 205.945 114.150 206.175 ;
        RECT 113.760 205.805 114.080 205.945 ;
        RECT 112.760 204.740 112.990 205.740 ;
        RECT 113.350 204.740 113.580 205.740 ;
        RECT 112.190 204.305 112.650 204.535 ;
        RECT 112.335 202.600 112.505 204.305 ;
        RECT 112.190 202.370 112.650 202.600 ;
        RECT 111.880 202.210 112.050 202.230 ;
        RECT 111.260 201.835 111.490 202.210 ;
        RECT 111.215 201.575 111.535 201.835 ;
        RECT 111.260 201.560 111.490 201.575 ;
        RECT 111.850 201.560 112.080 202.210 ;
        RECT 111.290 201.540 111.460 201.560 ;
        RECT 110.760 201.400 111.080 201.415 ;
        RECT 110.690 201.170 111.150 201.400 ;
        RECT 110.760 201.155 111.080 201.170 ;
        RECT 111.880 200.980 112.050 201.560 ;
        RECT 112.335 201.415 112.505 202.370 ;
        RECT 112.790 202.210 112.960 204.740 ;
        RECT 113.380 204.720 113.550 204.740 ;
        RECT 113.835 204.535 114.005 205.805 ;
        RECT 114.290 205.740 114.460 205.760 ;
        RECT 114.880 205.740 115.050 206.320 ;
        RECT 115.190 205.945 115.650 206.175 ;
        RECT 115.260 205.805 115.580 205.945 ;
        RECT 114.260 204.740 114.490 205.740 ;
        RECT 114.850 204.740 115.080 205.740 ;
        RECT 113.690 204.305 114.150 204.535 ;
        RECT 113.835 202.600 114.005 204.305 ;
        RECT 113.690 202.370 114.150 202.600 ;
        RECT 113.380 202.210 113.550 202.230 ;
        RECT 112.760 201.835 112.990 202.210 ;
        RECT 112.715 201.575 113.035 201.835 ;
        RECT 112.760 201.560 112.990 201.575 ;
        RECT 113.350 201.560 113.580 202.210 ;
        RECT 112.790 201.540 112.960 201.560 ;
        RECT 112.260 201.400 112.580 201.415 ;
        RECT 112.190 201.170 112.650 201.400 ;
        RECT 112.260 201.155 112.580 201.170 ;
        RECT 113.380 200.980 113.550 201.560 ;
        RECT 113.835 201.415 114.005 202.370 ;
        RECT 114.290 202.210 114.460 204.740 ;
        RECT 114.880 204.720 115.050 204.740 ;
        RECT 115.335 204.535 115.505 205.805 ;
        RECT 115.790 205.740 115.960 205.760 ;
        RECT 116.380 205.740 116.550 206.320 ;
        RECT 116.690 205.945 117.150 206.175 ;
        RECT 116.760 205.805 117.080 205.945 ;
        RECT 115.760 204.740 115.990 205.740 ;
        RECT 116.350 204.740 116.580 205.740 ;
        RECT 115.190 204.305 115.650 204.535 ;
        RECT 115.335 202.600 115.505 204.305 ;
        RECT 115.190 202.370 115.650 202.600 ;
        RECT 114.880 202.210 115.050 202.230 ;
        RECT 114.260 201.835 114.490 202.210 ;
        RECT 114.215 201.575 114.535 201.835 ;
        RECT 114.260 201.560 114.490 201.575 ;
        RECT 114.850 201.560 115.080 202.210 ;
        RECT 114.290 201.540 114.460 201.560 ;
        RECT 113.760 201.400 114.080 201.415 ;
        RECT 113.690 201.170 114.150 201.400 ;
        RECT 113.760 201.155 114.080 201.170 ;
        RECT 114.880 200.980 115.050 201.560 ;
        RECT 115.335 201.415 115.505 202.370 ;
        RECT 115.790 202.210 115.960 204.740 ;
        RECT 116.380 204.720 116.550 204.740 ;
        RECT 116.835 204.535 117.005 205.805 ;
        RECT 117.290 205.740 117.460 205.760 ;
        RECT 117.880 205.740 118.050 206.320 ;
        RECT 119.290 206.305 119.580 206.335 ;
        RECT 118.190 205.945 118.650 206.175 ;
        RECT 118.260 205.805 118.580 205.945 ;
        RECT 117.260 204.740 117.490 205.740 ;
        RECT 117.850 204.740 118.080 205.740 ;
        RECT 116.690 204.305 117.150 204.535 ;
        RECT 116.835 202.600 117.005 204.305 ;
        RECT 116.690 202.370 117.150 202.600 ;
        RECT 116.380 202.210 116.550 202.230 ;
        RECT 115.760 201.835 115.990 202.210 ;
        RECT 115.715 201.575 116.035 201.835 ;
        RECT 115.760 201.560 115.990 201.575 ;
        RECT 116.350 201.560 116.580 202.210 ;
        RECT 115.790 201.540 115.960 201.560 ;
        RECT 115.260 201.400 115.580 201.415 ;
        RECT 115.190 201.170 115.650 201.400 ;
        RECT 115.260 201.155 115.580 201.170 ;
        RECT 116.380 200.980 116.550 201.560 ;
        RECT 116.835 201.415 117.005 202.370 ;
        RECT 117.290 202.210 117.460 204.740 ;
        RECT 117.880 204.720 118.050 204.740 ;
        RECT 118.335 204.535 118.505 205.805 ;
        RECT 118.790 205.740 118.960 205.760 ;
        RECT 118.760 204.740 118.990 205.740 ;
        RECT 118.190 204.305 118.650 204.535 ;
        RECT 118.335 202.600 118.505 204.305 ;
        RECT 118.190 202.370 118.650 202.600 ;
        RECT 117.880 202.210 118.050 202.230 ;
        RECT 117.260 201.835 117.490 202.210 ;
        RECT 117.215 201.575 117.535 201.835 ;
        RECT 117.260 201.560 117.490 201.575 ;
        RECT 117.850 201.560 118.080 202.210 ;
        RECT 117.290 201.540 117.460 201.560 ;
        RECT 116.760 201.400 117.080 201.415 ;
        RECT 116.690 201.170 117.150 201.400 ;
        RECT 116.760 201.155 117.080 201.170 ;
        RECT 117.880 200.980 118.050 201.560 ;
        RECT 118.335 201.415 118.505 202.370 ;
        RECT 118.790 202.210 118.960 204.740 ;
        RECT 118.760 201.835 118.990 202.210 ;
        RECT 118.715 201.575 119.035 201.835 ;
        RECT 118.760 201.560 118.990 201.575 ;
        RECT 118.790 201.540 118.960 201.560 ;
        RECT 118.260 201.400 118.580 201.415 ;
        RECT 118.190 201.170 118.650 201.400 ;
        RECT 118.260 201.155 118.580 201.170 ;
        RECT 107.335 200.965 107.595 200.980 ;
        RECT 108.835 200.965 109.095 200.980 ;
        RECT 110.335 200.965 110.595 200.980 ;
        RECT 111.835 200.965 112.095 200.980 ;
        RECT 113.335 200.965 113.595 200.980 ;
        RECT 114.835 200.965 115.095 200.980 ;
        RECT 116.335 200.965 116.595 200.980 ;
        RECT 117.835 200.965 118.095 200.980 ;
        RECT 119.440 200.965 119.730 200.995 ;
        RECT 106.630 200.675 119.730 200.965 ;
        RECT 107.335 200.660 107.595 200.675 ;
        RECT 108.835 200.660 109.095 200.675 ;
        RECT 110.335 200.660 110.595 200.675 ;
        RECT 111.835 200.660 112.095 200.675 ;
        RECT 113.335 200.660 113.595 200.675 ;
        RECT 114.835 200.660 115.095 200.675 ;
        RECT 116.335 200.660 116.595 200.675 ;
        RECT 117.835 200.660 118.095 200.675 ;
        RECT 119.440 200.645 119.730 200.675 ;
        RECT 76.760 199.885 76.990 200.535 ;
        RECT 76.790 199.865 76.960 199.885 ;
        RECT 76.190 199.695 76.650 199.725 ;
        RECT 76.190 199.525 76.960 199.695 ;
        RECT 76.190 199.495 76.650 199.525 ;
        RECT 76.260 199.075 76.580 199.335 ;
        RECT 76.335 197.835 76.505 199.075 ;
        RECT 76.790 198.445 76.960 199.525 ;
        RECT 76.745 198.125 77.005 198.445 ;
        RECT 76.290 197.790 76.550 197.835 ;
        RECT 76.190 197.560 76.650 197.790 ;
        RECT 76.290 197.515 76.550 197.560 ;
        RECT 75.260 196.355 75.490 197.355 ;
        RECT 75.850 196.355 76.080 197.355 ;
        RECT 74.690 195.920 75.150 196.150 ;
        RECT 75.290 195.775 75.460 196.355 ;
        RECT 75.880 196.335 76.050 196.355 ;
        RECT 76.335 196.150 76.505 197.515 ;
        RECT 76.790 197.355 76.960 197.375 ;
        RECT 76.760 196.355 76.990 197.355 ;
        RECT 76.190 195.920 76.650 196.150 ;
        RECT 76.790 195.775 76.960 196.355 ;
        RECT 66.245 195.760 66.505 195.775 ;
        RECT 67.745 195.760 68.005 195.775 ;
        RECT 69.245 195.760 69.505 195.775 ;
        RECT 70.745 195.760 71.005 195.775 ;
        RECT 72.245 195.760 72.505 195.775 ;
        RECT 73.745 195.760 74.005 195.775 ;
        RECT 75.245 195.760 75.505 195.775 ;
        RECT 76.745 195.760 77.005 195.775 ;
        RECT 77.290 195.760 77.580 195.790 ;
        RECT 64.760 195.470 77.580 195.760 ;
        RECT 64.760 195.440 65.050 195.470 ;
        RECT 66.245 195.455 66.505 195.470 ;
        RECT 67.745 195.455 68.005 195.470 ;
        RECT 69.245 195.455 69.505 195.470 ;
        RECT 70.745 195.455 71.005 195.470 ;
        RECT 72.245 195.455 72.505 195.470 ;
        RECT 73.745 195.455 74.005 195.470 ;
        RECT 75.245 195.455 75.505 195.470 ;
        RECT 76.745 195.455 77.005 195.470 ;
        RECT 77.290 195.440 77.580 195.470 ;
        RECT 106.760 189.160 107.050 189.190 ;
        RECT 107.335 189.160 107.595 189.175 ;
        RECT 108.835 189.160 109.095 189.175 ;
        RECT 110.335 189.160 110.595 189.175 ;
        RECT 111.835 189.160 112.095 189.175 ;
        RECT 113.335 189.160 113.595 189.175 ;
        RECT 114.835 189.160 115.095 189.175 ;
        RECT 116.335 189.160 116.595 189.175 ;
        RECT 117.835 189.160 118.095 189.175 ;
        RECT 119.290 189.160 119.580 189.190 ;
        RECT 106.760 188.870 119.580 189.160 ;
        RECT 106.760 188.840 107.050 188.870 ;
        RECT 107.335 188.855 107.595 188.870 ;
        RECT 108.835 188.855 109.095 188.870 ;
        RECT 110.335 188.855 110.595 188.870 ;
        RECT 111.835 188.855 112.095 188.870 ;
        RECT 113.335 188.855 113.595 188.870 ;
        RECT 114.835 188.855 115.095 188.870 ;
        RECT 116.335 188.855 116.595 188.870 ;
        RECT 117.835 188.855 118.095 188.870 ;
        RECT 107.380 188.275 107.550 188.855 ;
        RECT 107.690 188.480 108.150 188.710 ;
        RECT 107.350 187.275 107.580 188.275 ;
        RECT 107.380 187.255 107.550 187.275 ;
        RECT 107.835 187.115 108.005 188.480 ;
        RECT 108.290 188.275 108.460 188.295 ;
        RECT 108.880 188.275 109.050 188.855 ;
        RECT 109.190 188.480 109.650 188.710 ;
        RECT 108.260 187.275 108.490 188.275 ;
        RECT 108.850 187.275 109.080 188.275 ;
        RECT 107.790 187.070 108.050 187.115 ;
        RECT 107.690 186.840 108.150 187.070 ;
        RECT 107.790 186.795 108.050 186.840 ;
        RECT 107.335 186.185 107.595 186.505 ;
        RECT 107.380 185.105 107.550 186.185 ;
        RECT 107.835 185.555 108.005 186.795 ;
        RECT 107.760 185.295 108.080 185.555 ;
        RECT 107.690 185.105 108.150 185.135 ;
        RECT 107.380 184.935 108.150 185.105 ;
        RECT 107.690 184.905 108.150 184.935 ;
        RECT 107.380 184.745 107.550 184.765 ;
        RECT 107.350 184.095 107.580 184.745 ;
        RECT 38.610 183.955 38.900 183.985 ;
        RECT 40.245 183.955 40.505 183.970 ;
        RECT 41.745 183.955 42.005 183.970 ;
        RECT 43.245 183.955 43.505 183.970 ;
        RECT 44.745 183.955 45.005 183.970 ;
        RECT 46.245 183.955 46.505 183.970 ;
        RECT 47.745 183.955 48.005 183.970 ;
        RECT 49.245 183.955 49.505 183.970 ;
        RECT 50.745 183.955 51.005 183.970 ;
        RECT 64.610 183.955 64.900 183.985 ;
        RECT 66.245 183.955 66.505 183.970 ;
        RECT 67.745 183.955 68.005 183.970 ;
        RECT 69.245 183.955 69.505 183.970 ;
        RECT 70.745 183.955 71.005 183.970 ;
        RECT 72.245 183.955 72.505 183.970 ;
        RECT 73.745 183.955 74.005 183.970 ;
        RECT 75.245 183.955 75.505 183.970 ;
        RECT 76.745 183.955 77.005 183.970 ;
        RECT 38.610 183.665 51.710 183.955 ;
        RECT 64.610 183.665 77.710 183.955 ;
        RECT 38.610 183.635 38.900 183.665 ;
        RECT 40.245 183.650 40.505 183.665 ;
        RECT 41.745 183.650 42.005 183.665 ;
        RECT 43.245 183.650 43.505 183.665 ;
        RECT 44.745 183.650 45.005 183.665 ;
        RECT 46.245 183.650 46.505 183.665 ;
        RECT 47.745 183.650 48.005 183.665 ;
        RECT 49.245 183.650 49.505 183.665 ;
        RECT 50.745 183.650 51.005 183.665 ;
        RECT 39.760 183.460 40.080 183.475 ;
        RECT 39.690 183.230 40.150 183.460 ;
        RECT 39.760 183.215 40.080 183.230 ;
        RECT 39.380 183.070 39.550 183.090 ;
        RECT 39.350 183.055 39.580 183.070 ;
        RECT 39.305 182.795 39.625 183.055 ;
        RECT 39.350 182.420 39.580 182.795 ;
        RECT 39.380 179.890 39.550 182.420 ;
        RECT 39.835 182.260 40.005 183.215 ;
        RECT 40.290 183.070 40.460 183.650 ;
        RECT 41.260 183.460 41.580 183.475 ;
        RECT 41.190 183.230 41.650 183.460 ;
        RECT 41.260 183.215 41.580 183.230 ;
        RECT 40.880 183.070 41.050 183.090 ;
        RECT 40.260 182.420 40.490 183.070 ;
        RECT 40.850 183.055 41.080 183.070 ;
        RECT 40.805 182.795 41.125 183.055 ;
        RECT 40.850 182.420 41.080 182.795 ;
        RECT 40.290 182.400 40.460 182.420 ;
        RECT 39.690 182.030 40.150 182.260 ;
        RECT 39.835 180.325 40.005 182.030 ;
        RECT 39.690 180.095 40.150 180.325 ;
        RECT 39.350 178.890 39.580 179.890 ;
        RECT 39.380 178.870 39.550 178.890 ;
        RECT 39.835 178.815 40.005 180.095 ;
        RECT 40.290 179.890 40.460 179.910 ;
        RECT 40.880 179.890 41.050 182.420 ;
        RECT 41.335 182.260 41.505 183.215 ;
        RECT 41.790 183.070 41.960 183.650 ;
        RECT 42.760 183.460 43.080 183.475 ;
        RECT 42.690 183.230 43.150 183.460 ;
        RECT 42.760 183.215 43.080 183.230 ;
        RECT 42.380 183.070 42.550 183.090 ;
        RECT 41.760 182.420 41.990 183.070 ;
        RECT 42.350 183.055 42.580 183.070 ;
        RECT 42.305 182.795 42.625 183.055 ;
        RECT 42.350 182.420 42.580 182.795 ;
        RECT 41.790 182.400 41.960 182.420 ;
        RECT 41.190 182.030 41.650 182.260 ;
        RECT 41.335 180.325 41.505 182.030 ;
        RECT 41.190 180.095 41.650 180.325 ;
        RECT 40.260 178.890 40.490 179.890 ;
        RECT 40.850 178.890 41.080 179.890 ;
        RECT 39.790 178.685 40.050 178.815 ;
        RECT 39.690 178.455 40.150 178.685 ;
        RECT 38.760 178.295 39.050 178.325 ;
        RECT 40.290 178.310 40.460 178.890 ;
        RECT 40.880 178.870 41.050 178.890 ;
        RECT 41.335 178.815 41.505 180.095 ;
        RECT 41.790 179.890 41.960 179.910 ;
        RECT 42.380 179.890 42.550 182.420 ;
        RECT 42.835 182.260 43.005 183.215 ;
        RECT 43.290 183.070 43.460 183.650 ;
        RECT 44.260 183.460 44.580 183.475 ;
        RECT 44.190 183.230 44.650 183.460 ;
        RECT 44.260 183.215 44.580 183.230 ;
        RECT 43.880 183.070 44.050 183.090 ;
        RECT 43.260 182.420 43.490 183.070 ;
        RECT 43.850 183.055 44.080 183.070 ;
        RECT 43.805 182.795 44.125 183.055 ;
        RECT 43.850 182.420 44.080 182.795 ;
        RECT 43.290 182.400 43.460 182.420 ;
        RECT 42.690 182.030 43.150 182.260 ;
        RECT 42.835 180.325 43.005 182.030 ;
        RECT 42.690 180.095 43.150 180.325 ;
        RECT 41.760 178.890 41.990 179.890 ;
        RECT 42.350 178.890 42.580 179.890 ;
        RECT 41.290 178.685 41.550 178.815 ;
        RECT 41.190 178.455 41.650 178.685 ;
        RECT 41.790 178.310 41.960 178.890 ;
        RECT 42.380 178.870 42.550 178.890 ;
        RECT 42.835 178.815 43.005 180.095 ;
        RECT 43.290 179.890 43.460 179.910 ;
        RECT 43.880 179.890 44.050 182.420 ;
        RECT 44.335 182.260 44.505 183.215 ;
        RECT 44.790 183.070 44.960 183.650 ;
        RECT 45.760 183.460 46.080 183.475 ;
        RECT 45.690 183.230 46.150 183.460 ;
        RECT 45.760 183.215 46.080 183.230 ;
        RECT 45.380 183.070 45.550 183.090 ;
        RECT 44.760 182.420 44.990 183.070 ;
        RECT 45.350 183.055 45.580 183.070 ;
        RECT 45.305 182.795 45.625 183.055 ;
        RECT 45.350 182.420 45.580 182.795 ;
        RECT 44.790 182.400 44.960 182.420 ;
        RECT 44.190 182.030 44.650 182.260 ;
        RECT 44.335 180.325 44.505 182.030 ;
        RECT 44.190 180.095 44.650 180.325 ;
        RECT 43.260 178.890 43.490 179.890 ;
        RECT 43.850 178.890 44.080 179.890 ;
        RECT 42.790 178.685 43.050 178.815 ;
        RECT 42.690 178.455 43.150 178.685 ;
        RECT 43.290 178.310 43.460 178.890 ;
        RECT 43.880 178.870 44.050 178.890 ;
        RECT 44.335 178.815 44.505 180.095 ;
        RECT 44.790 179.890 44.960 179.910 ;
        RECT 45.380 179.890 45.550 182.420 ;
        RECT 45.835 182.260 46.005 183.215 ;
        RECT 46.290 183.070 46.460 183.650 ;
        RECT 47.260 183.460 47.580 183.475 ;
        RECT 47.190 183.230 47.650 183.460 ;
        RECT 47.260 183.215 47.580 183.230 ;
        RECT 46.880 183.070 47.050 183.090 ;
        RECT 46.260 182.420 46.490 183.070 ;
        RECT 46.850 183.055 47.080 183.070 ;
        RECT 46.805 182.795 47.125 183.055 ;
        RECT 46.850 182.420 47.080 182.795 ;
        RECT 46.290 182.400 46.460 182.420 ;
        RECT 45.690 182.030 46.150 182.260 ;
        RECT 45.835 180.325 46.005 182.030 ;
        RECT 45.690 180.095 46.150 180.325 ;
        RECT 44.760 178.890 44.990 179.890 ;
        RECT 45.350 178.890 45.580 179.890 ;
        RECT 44.290 178.685 44.550 178.815 ;
        RECT 44.190 178.455 44.650 178.685 ;
        RECT 44.790 178.310 44.960 178.890 ;
        RECT 45.380 178.870 45.550 178.890 ;
        RECT 45.835 178.815 46.005 180.095 ;
        RECT 46.290 179.890 46.460 179.910 ;
        RECT 46.880 179.890 47.050 182.420 ;
        RECT 47.335 182.260 47.505 183.215 ;
        RECT 47.790 183.070 47.960 183.650 ;
        RECT 48.760 183.460 49.080 183.475 ;
        RECT 48.690 183.230 49.150 183.460 ;
        RECT 48.760 183.215 49.080 183.230 ;
        RECT 48.380 183.070 48.550 183.090 ;
        RECT 47.760 182.420 47.990 183.070 ;
        RECT 48.350 183.055 48.580 183.070 ;
        RECT 48.305 182.795 48.625 183.055 ;
        RECT 48.350 182.420 48.580 182.795 ;
        RECT 47.790 182.400 47.960 182.420 ;
        RECT 47.190 182.030 47.650 182.260 ;
        RECT 47.335 180.325 47.505 182.030 ;
        RECT 47.190 180.095 47.650 180.325 ;
        RECT 46.260 178.890 46.490 179.890 ;
        RECT 46.850 178.890 47.080 179.890 ;
        RECT 45.790 178.685 46.050 178.815 ;
        RECT 45.690 178.455 46.150 178.685 ;
        RECT 46.290 178.310 46.460 178.890 ;
        RECT 46.880 178.870 47.050 178.890 ;
        RECT 47.335 178.815 47.505 180.095 ;
        RECT 47.790 179.890 47.960 179.910 ;
        RECT 48.380 179.890 48.550 182.420 ;
        RECT 48.835 182.260 49.005 183.215 ;
        RECT 49.290 183.070 49.460 183.650 ;
        RECT 50.260 183.460 50.580 183.475 ;
        RECT 50.190 183.230 50.650 183.460 ;
        RECT 50.260 183.215 50.580 183.230 ;
        RECT 49.880 183.070 50.050 183.090 ;
        RECT 49.260 182.420 49.490 183.070 ;
        RECT 49.850 183.055 50.080 183.070 ;
        RECT 49.805 182.795 50.125 183.055 ;
        RECT 49.850 182.420 50.080 182.795 ;
        RECT 49.290 182.400 49.460 182.420 ;
        RECT 48.690 182.030 49.150 182.260 ;
        RECT 48.835 180.325 49.005 182.030 ;
        RECT 48.690 180.095 49.150 180.325 ;
        RECT 47.760 178.890 47.990 179.890 ;
        RECT 48.350 178.890 48.580 179.890 ;
        RECT 47.290 178.685 47.550 178.815 ;
        RECT 47.190 178.455 47.650 178.685 ;
        RECT 47.790 178.310 47.960 178.890 ;
        RECT 48.380 178.870 48.550 178.890 ;
        RECT 48.835 178.815 49.005 180.095 ;
        RECT 49.290 179.890 49.460 179.910 ;
        RECT 49.880 179.890 50.050 182.420 ;
        RECT 50.335 182.260 50.505 183.215 ;
        RECT 50.790 183.070 50.960 183.650 ;
        RECT 64.610 183.635 64.900 183.665 ;
        RECT 66.245 183.650 66.505 183.665 ;
        RECT 67.745 183.650 68.005 183.665 ;
        RECT 69.245 183.650 69.505 183.665 ;
        RECT 70.745 183.650 71.005 183.665 ;
        RECT 72.245 183.650 72.505 183.665 ;
        RECT 73.745 183.650 74.005 183.665 ;
        RECT 75.245 183.650 75.505 183.665 ;
        RECT 76.745 183.650 77.005 183.665 ;
        RECT 65.760 183.460 66.080 183.475 ;
        RECT 65.690 183.230 66.150 183.460 ;
        RECT 65.760 183.215 66.080 183.230 ;
        RECT 65.380 183.070 65.550 183.090 ;
        RECT 50.760 182.420 50.990 183.070 ;
        RECT 65.350 183.055 65.580 183.070 ;
        RECT 65.305 182.795 65.625 183.055 ;
        RECT 65.350 182.420 65.580 182.795 ;
        RECT 50.790 182.400 50.960 182.420 ;
        RECT 50.190 182.030 50.650 182.260 ;
        RECT 50.335 180.325 50.505 182.030 ;
        RECT 50.190 180.095 50.650 180.325 ;
        RECT 49.260 178.890 49.490 179.890 ;
        RECT 49.850 178.890 50.080 179.890 ;
        RECT 48.790 178.685 49.050 178.815 ;
        RECT 48.690 178.455 49.150 178.685 ;
        RECT 49.290 178.310 49.460 178.890 ;
        RECT 49.880 178.870 50.050 178.890 ;
        RECT 50.335 178.815 50.505 180.095 ;
        RECT 50.790 179.890 50.960 179.910 ;
        RECT 65.380 179.890 65.550 182.420 ;
        RECT 65.835 182.260 66.005 183.215 ;
        RECT 66.290 183.070 66.460 183.650 ;
        RECT 67.260 183.460 67.580 183.475 ;
        RECT 67.190 183.230 67.650 183.460 ;
        RECT 67.260 183.215 67.580 183.230 ;
        RECT 66.880 183.070 67.050 183.090 ;
        RECT 66.260 182.420 66.490 183.070 ;
        RECT 66.850 183.055 67.080 183.070 ;
        RECT 66.805 182.795 67.125 183.055 ;
        RECT 66.850 182.420 67.080 182.795 ;
        RECT 66.290 182.400 66.460 182.420 ;
        RECT 65.690 182.030 66.150 182.260 ;
        RECT 65.835 180.325 66.005 182.030 ;
        RECT 65.690 180.095 66.150 180.325 ;
        RECT 50.760 178.890 50.990 179.890 ;
        RECT 65.350 178.890 65.580 179.890 ;
        RECT 50.290 178.685 50.550 178.815 ;
        RECT 50.190 178.455 50.650 178.685 ;
        RECT 50.790 178.310 50.960 178.890 ;
        RECT 65.380 178.870 65.550 178.890 ;
        RECT 65.835 178.815 66.005 180.095 ;
        RECT 66.290 179.890 66.460 179.910 ;
        RECT 66.880 179.890 67.050 182.420 ;
        RECT 67.335 182.260 67.505 183.215 ;
        RECT 67.790 183.070 67.960 183.650 ;
        RECT 68.760 183.460 69.080 183.475 ;
        RECT 68.690 183.230 69.150 183.460 ;
        RECT 68.760 183.215 69.080 183.230 ;
        RECT 68.380 183.070 68.550 183.090 ;
        RECT 67.760 182.420 67.990 183.070 ;
        RECT 68.350 183.055 68.580 183.070 ;
        RECT 68.305 182.795 68.625 183.055 ;
        RECT 68.350 182.420 68.580 182.795 ;
        RECT 67.790 182.400 67.960 182.420 ;
        RECT 67.190 182.030 67.650 182.260 ;
        RECT 67.335 180.325 67.505 182.030 ;
        RECT 67.190 180.095 67.650 180.325 ;
        RECT 66.260 178.890 66.490 179.890 ;
        RECT 66.850 178.890 67.080 179.890 ;
        RECT 65.790 178.685 66.050 178.815 ;
        RECT 65.690 178.455 66.150 178.685 ;
        RECT 40.290 178.295 40.575 178.310 ;
        RECT 41.790 178.295 42.075 178.310 ;
        RECT 43.290 178.295 43.575 178.310 ;
        RECT 44.790 178.295 45.075 178.310 ;
        RECT 46.290 178.295 46.575 178.310 ;
        RECT 47.790 178.295 48.075 178.310 ;
        RECT 49.290 178.295 49.575 178.310 ;
        RECT 50.790 178.295 51.075 178.310 ;
        RECT 51.290 178.295 51.580 178.325 ;
        RECT 38.760 178.005 51.580 178.295 ;
        RECT 38.760 177.975 39.050 178.005 ;
        RECT 40.315 177.990 40.575 178.005 ;
        RECT 41.815 177.990 42.075 178.005 ;
        RECT 43.315 177.990 43.575 178.005 ;
        RECT 44.815 177.990 45.075 178.005 ;
        RECT 46.315 177.990 46.575 178.005 ;
        RECT 47.815 177.990 48.075 178.005 ;
        RECT 49.315 177.990 49.575 178.005 ;
        RECT 50.815 177.990 51.075 178.005 ;
        RECT 51.290 177.975 51.580 178.005 ;
        RECT 64.760 178.295 65.050 178.325 ;
        RECT 66.290 178.310 66.460 178.890 ;
        RECT 66.880 178.870 67.050 178.890 ;
        RECT 67.335 178.815 67.505 180.095 ;
        RECT 67.790 179.890 67.960 179.910 ;
        RECT 68.380 179.890 68.550 182.420 ;
        RECT 68.835 182.260 69.005 183.215 ;
        RECT 69.290 183.070 69.460 183.650 ;
        RECT 70.260 183.460 70.580 183.475 ;
        RECT 70.190 183.230 70.650 183.460 ;
        RECT 70.260 183.215 70.580 183.230 ;
        RECT 69.880 183.070 70.050 183.090 ;
        RECT 69.260 182.420 69.490 183.070 ;
        RECT 69.850 183.055 70.080 183.070 ;
        RECT 69.805 182.795 70.125 183.055 ;
        RECT 69.850 182.420 70.080 182.795 ;
        RECT 69.290 182.400 69.460 182.420 ;
        RECT 68.690 182.030 69.150 182.260 ;
        RECT 68.835 180.325 69.005 182.030 ;
        RECT 68.690 180.095 69.150 180.325 ;
        RECT 67.760 178.890 67.990 179.890 ;
        RECT 68.350 178.890 68.580 179.890 ;
        RECT 67.290 178.685 67.550 178.815 ;
        RECT 67.190 178.455 67.650 178.685 ;
        RECT 67.790 178.310 67.960 178.890 ;
        RECT 68.380 178.870 68.550 178.890 ;
        RECT 68.835 178.815 69.005 180.095 ;
        RECT 69.290 179.890 69.460 179.910 ;
        RECT 69.880 179.890 70.050 182.420 ;
        RECT 70.335 182.260 70.505 183.215 ;
        RECT 70.790 183.070 70.960 183.650 ;
        RECT 71.760 183.460 72.080 183.475 ;
        RECT 71.690 183.230 72.150 183.460 ;
        RECT 71.760 183.215 72.080 183.230 ;
        RECT 71.380 183.070 71.550 183.090 ;
        RECT 70.760 182.420 70.990 183.070 ;
        RECT 71.350 183.055 71.580 183.070 ;
        RECT 71.305 182.795 71.625 183.055 ;
        RECT 71.350 182.420 71.580 182.795 ;
        RECT 70.790 182.400 70.960 182.420 ;
        RECT 70.190 182.030 70.650 182.260 ;
        RECT 70.335 180.325 70.505 182.030 ;
        RECT 70.190 180.095 70.650 180.325 ;
        RECT 69.260 178.890 69.490 179.890 ;
        RECT 69.850 178.890 70.080 179.890 ;
        RECT 68.790 178.685 69.050 178.815 ;
        RECT 68.690 178.455 69.150 178.685 ;
        RECT 69.290 178.310 69.460 178.890 ;
        RECT 69.880 178.870 70.050 178.890 ;
        RECT 70.335 178.815 70.505 180.095 ;
        RECT 70.790 179.890 70.960 179.910 ;
        RECT 71.380 179.890 71.550 182.420 ;
        RECT 71.835 182.260 72.005 183.215 ;
        RECT 72.290 183.070 72.460 183.650 ;
        RECT 73.260 183.460 73.580 183.475 ;
        RECT 73.190 183.230 73.650 183.460 ;
        RECT 73.260 183.215 73.580 183.230 ;
        RECT 72.880 183.070 73.050 183.090 ;
        RECT 72.260 182.420 72.490 183.070 ;
        RECT 72.850 183.055 73.080 183.070 ;
        RECT 72.805 182.795 73.125 183.055 ;
        RECT 72.850 182.420 73.080 182.795 ;
        RECT 72.290 182.400 72.460 182.420 ;
        RECT 71.690 182.030 72.150 182.260 ;
        RECT 71.835 180.325 72.005 182.030 ;
        RECT 71.690 180.095 72.150 180.325 ;
        RECT 70.760 178.890 70.990 179.890 ;
        RECT 71.350 178.890 71.580 179.890 ;
        RECT 70.290 178.685 70.550 178.815 ;
        RECT 70.190 178.455 70.650 178.685 ;
        RECT 70.790 178.310 70.960 178.890 ;
        RECT 71.380 178.870 71.550 178.890 ;
        RECT 71.835 178.815 72.005 180.095 ;
        RECT 72.290 179.890 72.460 179.910 ;
        RECT 72.880 179.890 73.050 182.420 ;
        RECT 73.335 182.260 73.505 183.215 ;
        RECT 73.790 183.070 73.960 183.650 ;
        RECT 74.760 183.460 75.080 183.475 ;
        RECT 74.690 183.230 75.150 183.460 ;
        RECT 74.760 183.215 75.080 183.230 ;
        RECT 74.380 183.070 74.550 183.090 ;
        RECT 73.760 182.420 73.990 183.070 ;
        RECT 74.350 183.055 74.580 183.070 ;
        RECT 74.305 182.795 74.625 183.055 ;
        RECT 74.350 182.420 74.580 182.795 ;
        RECT 73.790 182.400 73.960 182.420 ;
        RECT 73.190 182.030 73.650 182.260 ;
        RECT 73.335 180.325 73.505 182.030 ;
        RECT 73.190 180.095 73.650 180.325 ;
        RECT 72.260 178.890 72.490 179.890 ;
        RECT 72.850 178.890 73.080 179.890 ;
        RECT 71.790 178.685 72.050 178.815 ;
        RECT 71.690 178.455 72.150 178.685 ;
        RECT 72.290 178.310 72.460 178.890 ;
        RECT 72.880 178.870 73.050 178.890 ;
        RECT 73.335 178.815 73.505 180.095 ;
        RECT 73.790 179.890 73.960 179.910 ;
        RECT 74.380 179.890 74.550 182.420 ;
        RECT 74.835 182.260 75.005 183.215 ;
        RECT 75.290 183.070 75.460 183.650 ;
        RECT 76.260 183.460 76.580 183.475 ;
        RECT 76.190 183.230 76.650 183.460 ;
        RECT 76.260 183.215 76.580 183.230 ;
        RECT 75.880 183.070 76.050 183.090 ;
        RECT 75.260 182.420 75.490 183.070 ;
        RECT 75.850 183.055 76.080 183.070 ;
        RECT 75.805 182.795 76.125 183.055 ;
        RECT 75.850 182.420 76.080 182.795 ;
        RECT 75.290 182.400 75.460 182.420 ;
        RECT 74.690 182.030 75.150 182.260 ;
        RECT 74.835 180.325 75.005 182.030 ;
        RECT 74.690 180.095 75.150 180.325 ;
        RECT 73.760 178.890 73.990 179.890 ;
        RECT 74.350 178.890 74.580 179.890 ;
        RECT 73.290 178.685 73.550 178.815 ;
        RECT 73.190 178.455 73.650 178.685 ;
        RECT 73.790 178.310 73.960 178.890 ;
        RECT 74.380 178.870 74.550 178.890 ;
        RECT 74.835 178.815 75.005 180.095 ;
        RECT 75.290 179.890 75.460 179.910 ;
        RECT 75.880 179.890 76.050 182.420 ;
        RECT 76.335 182.260 76.505 183.215 ;
        RECT 76.790 183.070 76.960 183.650 ;
        RECT 106.630 183.500 106.980 183.560 ;
        RECT 107.380 183.500 107.550 184.095 ;
        RECT 107.835 183.935 108.005 184.905 ;
        RECT 108.290 184.745 108.460 187.275 ;
        RECT 108.880 187.255 109.050 187.275 ;
        RECT 109.335 187.115 109.505 188.480 ;
        RECT 109.790 188.275 109.960 188.295 ;
        RECT 110.380 188.275 110.550 188.855 ;
        RECT 110.690 188.480 111.150 188.710 ;
        RECT 109.760 187.275 109.990 188.275 ;
        RECT 110.350 187.275 110.580 188.275 ;
        RECT 109.290 187.070 109.550 187.115 ;
        RECT 109.190 186.840 109.650 187.070 ;
        RECT 109.290 186.795 109.550 186.840 ;
        RECT 108.835 186.185 109.095 186.505 ;
        RECT 108.880 185.105 109.050 186.185 ;
        RECT 109.335 185.555 109.505 186.795 ;
        RECT 109.260 185.295 109.580 185.555 ;
        RECT 109.190 185.105 109.650 185.135 ;
        RECT 108.880 184.935 109.650 185.105 ;
        RECT 109.190 184.905 109.650 184.935 ;
        RECT 108.880 184.745 109.050 184.765 ;
        RECT 108.260 184.400 108.490 184.745 ;
        RECT 108.245 184.080 108.505 184.400 ;
        RECT 108.850 184.095 109.080 184.745 ;
        RECT 108.290 184.075 108.460 184.080 ;
        RECT 107.690 183.705 108.150 183.935 ;
        RECT 108.880 183.500 109.050 184.095 ;
        RECT 109.335 183.935 109.505 184.905 ;
        RECT 109.790 184.745 109.960 187.275 ;
        RECT 110.380 187.255 110.550 187.275 ;
        RECT 110.835 187.115 111.005 188.480 ;
        RECT 111.290 188.275 111.460 188.295 ;
        RECT 111.880 188.275 112.050 188.855 ;
        RECT 112.190 188.480 112.650 188.710 ;
        RECT 111.260 187.275 111.490 188.275 ;
        RECT 111.850 187.275 112.080 188.275 ;
        RECT 110.790 187.070 111.050 187.115 ;
        RECT 110.690 186.840 111.150 187.070 ;
        RECT 110.790 186.795 111.050 186.840 ;
        RECT 110.335 186.185 110.595 186.505 ;
        RECT 110.380 185.105 110.550 186.185 ;
        RECT 110.835 185.555 111.005 186.795 ;
        RECT 110.760 185.295 111.080 185.555 ;
        RECT 110.690 185.105 111.150 185.135 ;
        RECT 110.380 184.935 111.150 185.105 ;
        RECT 110.690 184.905 111.150 184.935 ;
        RECT 110.380 184.745 110.550 184.765 ;
        RECT 109.760 184.400 109.990 184.745 ;
        RECT 109.745 184.080 110.005 184.400 ;
        RECT 110.350 184.095 110.580 184.745 ;
        RECT 109.790 184.075 109.960 184.080 ;
        RECT 109.190 183.705 109.650 183.935 ;
        RECT 110.380 183.500 110.550 184.095 ;
        RECT 110.835 183.935 111.005 184.905 ;
        RECT 111.290 184.745 111.460 187.275 ;
        RECT 111.880 187.255 112.050 187.275 ;
        RECT 112.335 187.115 112.505 188.480 ;
        RECT 112.790 188.275 112.960 188.295 ;
        RECT 113.380 188.275 113.550 188.855 ;
        RECT 113.690 188.480 114.150 188.710 ;
        RECT 112.760 187.275 112.990 188.275 ;
        RECT 113.350 187.275 113.580 188.275 ;
        RECT 112.290 187.070 112.550 187.115 ;
        RECT 112.190 186.840 112.650 187.070 ;
        RECT 112.290 186.795 112.550 186.840 ;
        RECT 111.835 186.185 112.095 186.505 ;
        RECT 111.880 185.105 112.050 186.185 ;
        RECT 112.335 185.555 112.505 186.795 ;
        RECT 112.260 185.295 112.580 185.555 ;
        RECT 112.190 185.105 112.650 185.135 ;
        RECT 111.880 184.935 112.650 185.105 ;
        RECT 112.190 184.905 112.650 184.935 ;
        RECT 111.880 184.745 112.050 184.765 ;
        RECT 111.260 184.400 111.490 184.745 ;
        RECT 111.245 184.080 111.505 184.400 ;
        RECT 111.850 184.095 112.080 184.745 ;
        RECT 111.290 184.075 111.460 184.080 ;
        RECT 110.690 183.705 111.150 183.935 ;
        RECT 111.880 183.500 112.050 184.095 ;
        RECT 112.335 183.935 112.505 184.905 ;
        RECT 112.790 184.745 112.960 187.275 ;
        RECT 113.380 187.255 113.550 187.275 ;
        RECT 113.835 187.115 114.005 188.480 ;
        RECT 114.290 188.275 114.460 188.295 ;
        RECT 114.880 188.275 115.050 188.855 ;
        RECT 115.190 188.480 115.650 188.710 ;
        RECT 114.260 187.275 114.490 188.275 ;
        RECT 114.850 187.275 115.080 188.275 ;
        RECT 113.790 187.070 114.050 187.115 ;
        RECT 113.690 186.840 114.150 187.070 ;
        RECT 113.790 186.795 114.050 186.840 ;
        RECT 113.335 186.185 113.595 186.505 ;
        RECT 113.380 185.105 113.550 186.185 ;
        RECT 113.835 185.555 114.005 186.795 ;
        RECT 113.760 185.295 114.080 185.555 ;
        RECT 113.690 185.105 114.150 185.135 ;
        RECT 113.380 184.935 114.150 185.105 ;
        RECT 113.690 184.905 114.150 184.935 ;
        RECT 113.380 184.745 113.550 184.765 ;
        RECT 112.760 184.400 112.990 184.745 ;
        RECT 112.745 184.080 113.005 184.400 ;
        RECT 113.350 184.095 113.580 184.745 ;
        RECT 112.790 184.075 112.960 184.080 ;
        RECT 112.190 183.705 112.650 183.935 ;
        RECT 113.380 183.500 113.550 184.095 ;
        RECT 113.835 183.935 114.005 184.905 ;
        RECT 114.290 184.745 114.460 187.275 ;
        RECT 114.880 187.255 115.050 187.275 ;
        RECT 115.335 187.115 115.505 188.480 ;
        RECT 115.790 188.275 115.960 188.295 ;
        RECT 116.380 188.275 116.550 188.855 ;
        RECT 116.690 188.480 117.150 188.710 ;
        RECT 115.760 187.275 115.990 188.275 ;
        RECT 116.350 187.275 116.580 188.275 ;
        RECT 115.290 187.070 115.550 187.115 ;
        RECT 115.190 186.840 115.650 187.070 ;
        RECT 115.290 186.795 115.550 186.840 ;
        RECT 114.835 186.185 115.095 186.505 ;
        RECT 114.880 185.105 115.050 186.185 ;
        RECT 115.335 185.555 115.505 186.795 ;
        RECT 115.260 185.295 115.580 185.555 ;
        RECT 115.190 185.105 115.650 185.135 ;
        RECT 114.880 184.935 115.650 185.105 ;
        RECT 115.190 184.905 115.650 184.935 ;
        RECT 114.880 184.745 115.050 184.765 ;
        RECT 114.260 184.400 114.490 184.745 ;
        RECT 114.245 184.080 114.505 184.400 ;
        RECT 114.850 184.095 115.080 184.745 ;
        RECT 114.290 184.075 114.460 184.080 ;
        RECT 113.690 183.705 114.150 183.935 ;
        RECT 114.880 183.500 115.050 184.095 ;
        RECT 115.335 183.935 115.505 184.905 ;
        RECT 115.790 184.745 115.960 187.275 ;
        RECT 116.380 187.255 116.550 187.275 ;
        RECT 116.835 187.115 117.005 188.480 ;
        RECT 117.290 188.275 117.460 188.295 ;
        RECT 117.880 188.275 118.050 188.855 ;
        RECT 119.290 188.840 119.580 188.870 ;
        RECT 118.190 188.480 118.650 188.710 ;
        RECT 117.260 187.275 117.490 188.275 ;
        RECT 117.850 187.275 118.080 188.275 ;
        RECT 116.790 187.070 117.050 187.115 ;
        RECT 116.690 186.840 117.150 187.070 ;
        RECT 116.790 186.795 117.050 186.840 ;
        RECT 116.335 186.185 116.595 186.505 ;
        RECT 116.380 185.105 116.550 186.185 ;
        RECT 116.835 185.555 117.005 186.795 ;
        RECT 116.760 185.295 117.080 185.555 ;
        RECT 116.690 185.105 117.150 185.135 ;
        RECT 116.380 184.935 117.150 185.105 ;
        RECT 116.690 184.905 117.150 184.935 ;
        RECT 116.380 184.745 116.550 184.765 ;
        RECT 115.760 184.400 115.990 184.745 ;
        RECT 115.745 184.080 116.005 184.400 ;
        RECT 116.350 184.095 116.580 184.745 ;
        RECT 115.790 184.075 115.960 184.080 ;
        RECT 115.190 183.705 115.650 183.935 ;
        RECT 116.380 183.500 116.550 184.095 ;
        RECT 116.835 183.935 117.005 184.905 ;
        RECT 117.290 184.745 117.460 187.275 ;
        RECT 117.880 187.255 118.050 187.275 ;
        RECT 118.335 187.115 118.505 188.480 ;
        RECT 118.790 188.275 118.960 188.295 ;
        RECT 118.760 187.275 118.990 188.275 ;
        RECT 118.290 187.070 118.550 187.115 ;
        RECT 118.190 186.840 118.650 187.070 ;
        RECT 118.290 186.795 118.550 186.840 ;
        RECT 117.835 186.185 118.095 186.505 ;
        RECT 117.880 185.105 118.050 186.185 ;
        RECT 118.335 185.555 118.505 186.795 ;
        RECT 118.260 185.295 118.580 185.555 ;
        RECT 118.190 185.105 118.650 185.135 ;
        RECT 117.880 184.935 118.650 185.105 ;
        RECT 118.190 184.905 118.650 184.935 ;
        RECT 117.880 184.745 118.050 184.765 ;
        RECT 117.260 184.400 117.490 184.745 ;
        RECT 117.245 184.080 117.505 184.400 ;
        RECT 117.850 184.095 118.080 184.745 ;
        RECT 117.290 184.075 117.460 184.080 ;
        RECT 116.690 183.705 117.150 183.935 ;
        RECT 117.880 183.500 118.050 184.095 ;
        RECT 118.335 183.935 118.505 184.905 ;
        RECT 118.790 184.745 118.960 187.275 ;
        RECT 118.760 184.400 118.990 184.745 ;
        RECT 118.745 184.080 119.005 184.400 ;
        RECT 118.790 184.075 118.960 184.080 ;
        RECT 118.190 183.705 118.650 183.935 ;
        RECT 119.410 183.500 119.760 183.560 ;
        RECT 106.630 183.210 119.760 183.500 ;
        RECT 106.630 183.150 106.980 183.210 ;
        RECT 119.410 183.150 119.760 183.210 ;
        RECT 76.760 182.420 76.990 183.070 ;
        RECT 106.730 182.450 107.080 182.510 ;
        RECT 119.265 182.450 119.615 182.510 ;
        RECT 76.790 182.400 76.960 182.420 ;
        RECT 76.190 182.030 76.650 182.260 ;
        RECT 106.730 182.160 119.615 182.450 ;
        RECT 106.730 182.100 107.080 182.160 ;
        RECT 76.335 180.325 76.505 182.030 ;
        RECT 107.380 181.565 107.550 182.160 ;
        RECT 107.690 181.970 108.150 182.000 ;
        RECT 108.310 181.970 108.630 182.015 ;
        RECT 107.690 181.800 108.630 181.970 ;
        RECT 107.690 181.770 108.150 181.800 ;
        RECT 107.350 180.565 107.580 181.565 ;
        RECT 107.380 180.545 107.550 180.565 ;
        RECT 107.835 180.360 108.005 181.770 ;
        RECT 108.310 181.755 108.630 181.800 ;
        RECT 108.290 181.565 108.460 181.585 ;
        RECT 108.880 181.565 109.050 182.160 ;
        RECT 109.190 181.970 109.650 182.000 ;
        RECT 109.810 181.970 110.130 182.015 ;
        RECT 109.190 181.800 110.130 181.970 ;
        RECT 109.190 181.770 109.650 181.800 ;
        RECT 108.260 181.530 108.490 181.565 ;
        RECT 108.215 181.270 108.535 181.530 ;
        RECT 108.260 180.565 108.490 181.270 ;
        RECT 108.850 180.565 109.080 181.565 ;
        RECT 76.190 180.095 76.650 180.325 ;
        RECT 107.690 180.130 108.150 180.360 ;
        RECT 75.260 178.890 75.490 179.890 ;
        RECT 75.850 178.890 76.080 179.890 ;
        RECT 74.790 178.685 75.050 178.815 ;
        RECT 74.690 178.455 75.150 178.685 ;
        RECT 75.290 178.310 75.460 178.890 ;
        RECT 75.880 178.870 76.050 178.890 ;
        RECT 76.335 178.815 76.505 180.095 ;
        RECT 76.790 179.890 76.960 179.910 ;
        RECT 76.760 178.890 76.990 179.890 ;
        RECT 76.290 178.685 76.550 178.815 ;
        RECT 76.190 178.455 76.650 178.685 ;
        RECT 76.790 178.310 76.960 178.890 ;
        RECT 107.790 178.425 108.050 178.470 ;
        RECT 66.290 178.295 66.575 178.310 ;
        RECT 67.790 178.295 68.075 178.310 ;
        RECT 69.290 178.295 69.575 178.310 ;
        RECT 70.790 178.295 71.075 178.310 ;
        RECT 72.290 178.295 72.575 178.310 ;
        RECT 73.790 178.295 74.075 178.310 ;
        RECT 75.290 178.295 75.575 178.310 ;
        RECT 76.790 178.295 77.075 178.310 ;
        RECT 77.290 178.295 77.580 178.325 ;
        RECT 64.760 178.005 77.580 178.295 ;
        RECT 107.690 178.195 108.150 178.425 ;
        RECT 107.790 178.150 108.050 178.195 ;
        RECT 107.380 178.035 107.550 178.055 ;
        RECT 64.760 177.975 65.050 178.005 ;
        RECT 66.315 177.990 66.575 178.005 ;
        RECT 67.815 177.990 68.075 178.005 ;
        RECT 69.315 177.990 69.575 178.005 ;
        RECT 70.815 177.990 71.075 178.005 ;
        RECT 72.315 177.990 72.575 178.005 ;
        RECT 73.815 177.990 74.075 178.005 ;
        RECT 75.315 177.990 75.575 178.005 ;
        RECT 76.815 177.990 77.075 178.005 ;
        RECT 77.290 177.975 77.580 178.005 ;
        RECT 107.350 177.385 107.580 178.035 ;
        RECT 106.660 176.790 106.950 176.820 ;
        RECT 107.380 176.805 107.550 177.385 ;
        RECT 107.835 177.225 108.005 178.150 ;
        RECT 108.290 178.035 108.460 180.565 ;
        RECT 108.880 180.545 109.050 180.565 ;
        RECT 109.335 180.360 109.505 181.770 ;
        RECT 109.810 181.755 110.130 181.800 ;
        RECT 109.790 181.565 109.960 181.585 ;
        RECT 110.380 181.565 110.550 182.160 ;
        RECT 110.690 181.970 111.150 182.000 ;
        RECT 111.310 181.970 111.630 182.015 ;
        RECT 110.690 181.800 111.630 181.970 ;
        RECT 110.690 181.770 111.150 181.800 ;
        RECT 109.760 181.530 109.990 181.565 ;
        RECT 109.715 181.270 110.035 181.530 ;
        RECT 109.760 180.565 109.990 181.270 ;
        RECT 110.350 180.565 110.580 181.565 ;
        RECT 109.190 180.130 109.650 180.360 ;
        RECT 109.290 178.425 109.550 178.470 ;
        RECT 109.190 178.195 109.650 178.425 ;
        RECT 109.290 178.150 109.550 178.195 ;
        RECT 108.880 178.035 109.050 178.055 ;
        RECT 108.260 177.690 108.490 178.035 ;
        RECT 108.245 177.370 108.505 177.690 ;
        RECT 108.850 177.385 109.080 178.035 ;
        RECT 108.290 177.365 108.460 177.370 ;
        RECT 107.690 176.995 108.150 177.225 ;
        RECT 108.880 176.805 109.050 177.385 ;
        RECT 109.335 177.225 109.505 178.150 ;
        RECT 109.790 178.035 109.960 180.565 ;
        RECT 110.380 180.545 110.550 180.565 ;
        RECT 110.835 180.360 111.005 181.770 ;
        RECT 111.310 181.755 111.630 181.800 ;
        RECT 111.290 181.565 111.460 181.585 ;
        RECT 111.880 181.565 112.050 182.160 ;
        RECT 112.190 181.970 112.650 182.000 ;
        RECT 112.810 181.970 113.130 182.015 ;
        RECT 112.190 181.800 113.130 181.970 ;
        RECT 112.190 181.770 112.650 181.800 ;
        RECT 111.260 181.530 111.490 181.565 ;
        RECT 111.215 181.270 111.535 181.530 ;
        RECT 111.260 180.565 111.490 181.270 ;
        RECT 111.850 180.565 112.080 181.565 ;
        RECT 110.690 180.130 111.150 180.360 ;
        RECT 110.790 178.425 111.050 178.470 ;
        RECT 110.690 178.195 111.150 178.425 ;
        RECT 110.790 178.150 111.050 178.195 ;
        RECT 110.380 178.035 110.550 178.055 ;
        RECT 109.760 177.690 109.990 178.035 ;
        RECT 109.745 177.370 110.005 177.690 ;
        RECT 110.350 177.385 110.580 178.035 ;
        RECT 109.790 177.365 109.960 177.370 ;
        RECT 109.190 176.995 109.650 177.225 ;
        RECT 110.380 176.805 110.550 177.385 ;
        RECT 110.835 177.225 111.005 178.150 ;
        RECT 111.290 178.035 111.460 180.565 ;
        RECT 111.880 180.545 112.050 180.565 ;
        RECT 112.335 180.360 112.505 181.770 ;
        RECT 112.810 181.755 113.130 181.800 ;
        RECT 112.790 181.565 112.960 181.585 ;
        RECT 113.380 181.565 113.550 182.160 ;
        RECT 113.690 181.970 114.150 182.000 ;
        RECT 114.310 181.970 114.630 182.015 ;
        RECT 113.690 181.800 114.630 181.970 ;
        RECT 113.690 181.770 114.150 181.800 ;
        RECT 112.760 181.530 112.990 181.565 ;
        RECT 112.715 181.270 113.035 181.530 ;
        RECT 112.760 180.565 112.990 181.270 ;
        RECT 113.350 180.565 113.580 181.565 ;
        RECT 112.190 180.130 112.650 180.360 ;
        RECT 112.290 178.425 112.550 178.470 ;
        RECT 112.190 178.195 112.650 178.425 ;
        RECT 112.290 178.150 112.550 178.195 ;
        RECT 111.880 178.035 112.050 178.055 ;
        RECT 111.260 177.690 111.490 178.035 ;
        RECT 111.245 177.370 111.505 177.690 ;
        RECT 111.850 177.385 112.080 178.035 ;
        RECT 111.290 177.365 111.460 177.370 ;
        RECT 110.690 176.995 111.150 177.225 ;
        RECT 111.880 176.805 112.050 177.385 ;
        RECT 112.335 177.225 112.505 178.150 ;
        RECT 112.790 178.035 112.960 180.565 ;
        RECT 113.380 180.545 113.550 180.565 ;
        RECT 113.835 180.360 114.005 181.770 ;
        RECT 114.310 181.755 114.630 181.800 ;
        RECT 114.290 181.565 114.460 181.585 ;
        RECT 114.880 181.565 115.050 182.160 ;
        RECT 115.190 181.970 115.650 182.000 ;
        RECT 115.810 181.970 116.130 182.015 ;
        RECT 115.190 181.800 116.130 181.970 ;
        RECT 115.190 181.770 115.650 181.800 ;
        RECT 114.260 181.530 114.490 181.565 ;
        RECT 114.215 181.270 114.535 181.530 ;
        RECT 114.260 180.565 114.490 181.270 ;
        RECT 114.850 180.565 115.080 181.565 ;
        RECT 113.690 180.130 114.150 180.360 ;
        RECT 113.790 178.425 114.050 178.470 ;
        RECT 113.690 178.195 114.150 178.425 ;
        RECT 113.790 178.150 114.050 178.195 ;
        RECT 113.380 178.035 113.550 178.055 ;
        RECT 112.760 177.690 112.990 178.035 ;
        RECT 112.745 177.370 113.005 177.690 ;
        RECT 113.350 177.385 113.580 178.035 ;
        RECT 112.790 177.365 112.960 177.370 ;
        RECT 112.190 176.995 112.650 177.225 ;
        RECT 113.380 176.805 113.550 177.385 ;
        RECT 113.835 177.225 114.005 178.150 ;
        RECT 114.290 178.035 114.460 180.565 ;
        RECT 114.880 180.545 115.050 180.565 ;
        RECT 115.335 180.360 115.505 181.770 ;
        RECT 115.810 181.755 116.130 181.800 ;
        RECT 115.790 181.565 115.960 181.585 ;
        RECT 116.380 181.565 116.550 182.160 ;
        RECT 116.690 181.970 117.150 182.000 ;
        RECT 117.310 181.970 117.630 182.015 ;
        RECT 116.690 181.800 117.630 181.970 ;
        RECT 116.690 181.770 117.150 181.800 ;
        RECT 115.760 181.530 115.990 181.565 ;
        RECT 115.715 181.270 116.035 181.530 ;
        RECT 115.760 180.565 115.990 181.270 ;
        RECT 116.350 180.565 116.580 181.565 ;
        RECT 115.190 180.130 115.650 180.360 ;
        RECT 115.290 178.425 115.550 178.470 ;
        RECT 115.190 178.195 115.650 178.425 ;
        RECT 115.290 178.150 115.550 178.195 ;
        RECT 114.880 178.035 115.050 178.055 ;
        RECT 114.260 177.690 114.490 178.035 ;
        RECT 114.245 177.370 114.505 177.690 ;
        RECT 114.850 177.385 115.080 178.035 ;
        RECT 114.290 177.365 114.460 177.370 ;
        RECT 113.690 176.995 114.150 177.225 ;
        RECT 114.880 176.805 115.050 177.385 ;
        RECT 115.335 177.225 115.505 178.150 ;
        RECT 115.790 178.035 115.960 180.565 ;
        RECT 116.380 180.545 116.550 180.565 ;
        RECT 116.835 180.360 117.005 181.770 ;
        RECT 117.310 181.755 117.630 181.800 ;
        RECT 117.290 181.565 117.460 181.585 ;
        RECT 117.880 181.565 118.050 182.160 ;
        RECT 119.265 182.100 119.615 182.160 ;
        RECT 118.190 181.970 118.650 182.000 ;
        RECT 118.810 181.970 119.130 182.015 ;
        RECT 118.190 181.800 119.130 181.970 ;
        RECT 118.190 181.770 118.650 181.800 ;
        RECT 117.260 181.530 117.490 181.565 ;
        RECT 117.215 181.270 117.535 181.530 ;
        RECT 117.260 180.565 117.490 181.270 ;
        RECT 117.850 180.565 118.080 181.565 ;
        RECT 116.690 180.130 117.150 180.360 ;
        RECT 116.790 178.425 117.050 178.470 ;
        RECT 116.690 178.195 117.150 178.425 ;
        RECT 116.790 178.150 117.050 178.195 ;
        RECT 116.380 178.035 116.550 178.055 ;
        RECT 115.760 177.690 115.990 178.035 ;
        RECT 115.745 177.370 116.005 177.690 ;
        RECT 116.350 177.385 116.580 178.035 ;
        RECT 115.790 177.365 115.960 177.370 ;
        RECT 115.190 176.995 115.650 177.225 ;
        RECT 116.380 176.805 116.550 177.385 ;
        RECT 116.835 177.225 117.005 178.150 ;
        RECT 117.290 178.035 117.460 180.565 ;
        RECT 117.880 180.545 118.050 180.565 ;
        RECT 118.335 180.360 118.505 181.770 ;
        RECT 118.810 181.755 119.130 181.800 ;
        RECT 118.790 181.565 118.960 181.585 ;
        RECT 118.760 181.530 118.990 181.565 ;
        RECT 118.715 181.270 119.035 181.530 ;
        RECT 118.760 180.565 118.990 181.270 ;
        RECT 118.190 180.130 118.650 180.360 ;
        RECT 118.290 178.425 118.550 178.470 ;
        RECT 118.190 178.195 118.650 178.425 ;
        RECT 118.290 178.150 118.550 178.195 ;
        RECT 117.880 178.035 118.050 178.055 ;
        RECT 117.260 177.690 117.490 178.035 ;
        RECT 117.245 177.370 117.505 177.690 ;
        RECT 117.850 177.385 118.080 178.035 ;
        RECT 117.290 177.365 117.460 177.370 ;
        RECT 116.690 176.995 117.150 177.225 ;
        RECT 117.880 176.805 118.050 177.385 ;
        RECT 118.335 177.225 118.505 178.150 ;
        RECT 118.790 178.035 118.960 180.565 ;
        RECT 118.760 177.690 118.990 178.035 ;
        RECT 118.745 177.370 119.005 177.690 ;
        RECT 118.790 177.365 118.960 177.370 ;
        RECT 118.190 176.995 118.650 177.225 ;
        RECT 107.330 176.790 107.590 176.805 ;
        RECT 108.830 176.790 109.090 176.805 ;
        RECT 110.330 176.790 110.590 176.805 ;
        RECT 111.830 176.790 112.090 176.805 ;
        RECT 113.330 176.790 113.590 176.805 ;
        RECT 114.830 176.790 115.090 176.805 ;
        RECT 116.330 176.790 116.590 176.805 ;
        RECT 117.830 176.790 118.090 176.805 ;
        RECT 119.440 176.790 119.730 176.820 ;
        RECT 106.660 176.500 119.730 176.790 ;
        RECT 106.660 176.470 106.950 176.500 ;
        RECT 107.330 176.485 107.590 176.500 ;
        RECT 108.830 176.485 109.090 176.500 ;
        RECT 110.330 176.485 110.590 176.500 ;
        RECT 111.830 176.485 112.090 176.500 ;
        RECT 113.330 176.485 113.590 176.500 ;
        RECT 114.830 176.485 115.090 176.500 ;
        RECT 116.330 176.485 116.590 176.500 ;
        RECT 117.830 176.485 118.090 176.500 ;
        RECT 119.440 176.470 119.730 176.500 ;
        RECT 38.595 167.845 38.945 167.875 ;
        RECT 43.155 167.845 43.505 167.875 ;
        RECT 38.595 167.495 43.505 167.845 ;
        RECT 38.595 167.465 38.945 167.495 ;
        RECT 43.155 167.465 43.505 167.495 ;
        RECT 40.875 166.845 41.225 166.875 ;
        RECT 69.995 166.845 70.345 166.875 ;
        RECT 40.875 166.495 70.345 166.845 ;
        RECT 40.875 166.465 41.225 166.495 ;
        RECT 69.995 166.465 70.345 166.495 ;
        RECT 39.670 165.845 40.020 165.875 ;
        RECT 41.950 165.845 42.300 165.875 ;
        RECT 39.670 165.495 42.300 165.845 ;
        RECT 39.670 165.465 40.020 165.495 ;
        RECT 41.950 165.465 42.300 165.495 ;
        RECT 44.230 164.845 44.580 164.875 ;
        RECT 66.510 164.845 66.860 164.875 ;
        RECT 44.230 164.495 66.860 164.845 ;
        RECT 44.230 164.465 44.580 164.495 ;
        RECT 66.510 164.465 66.860 164.495 ;
        RECT 45.305 163.845 45.655 163.875 ;
        RECT 49.865 163.845 50.215 163.875 ;
        RECT 45.305 163.495 50.215 163.845 ;
        RECT 45.305 163.465 45.655 163.495 ;
        RECT 49.865 163.465 50.215 163.495 ;
        RECT 47.585 162.845 47.935 162.875 ;
        RECT 76.705 162.845 77.055 162.875 ;
        RECT 47.585 162.495 77.055 162.845 ;
        RECT 47.585 162.465 47.935 162.495 ;
        RECT 76.705 162.465 77.055 162.495 ;
        RECT 46.380 161.845 46.730 161.875 ;
        RECT 48.660 161.845 49.010 161.875 ;
        RECT 46.380 161.495 49.010 161.845 ;
        RECT 46.380 161.465 46.730 161.495 ;
        RECT 48.660 161.465 49.010 161.495 ;
        RECT 50.940 160.845 51.290 160.875 ;
        RECT 73.220 160.845 73.570 160.875 ;
        RECT 50.940 160.495 73.570 160.845 ;
        RECT 50.940 160.465 51.290 160.495 ;
        RECT 73.220 160.465 73.570 160.495 ;
        RECT 29.735 159.845 30.085 159.875 ;
        RECT 65.435 159.845 65.785 159.875 ;
        RECT 29.735 159.495 65.785 159.845 ;
        RECT 29.735 159.465 30.085 159.495 ;
        RECT 65.435 159.465 65.785 159.495 ;
        RECT 56.575 158.845 56.925 158.875 ;
        RECT 67.715 158.845 68.065 158.875 ;
        RECT 56.575 158.495 68.065 158.845 ;
        RECT 56.575 158.465 56.925 158.495 ;
        RECT 67.715 158.465 68.065 158.495 ;
        RECT 26.250 157.845 26.600 157.875 ;
        RECT 68.790 157.845 69.140 157.875 ;
        RECT 26.250 157.495 69.140 157.845 ;
        RECT 26.250 157.465 26.600 157.495 ;
        RECT 68.790 157.465 69.140 157.495 ;
        RECT 53.090 156.845 53.440 156.875 ;
        RECT 71.070 156.845 71.420 156.875 ;
        RECT 53.090 156.495 71.420 156.845 ;
        RECT 53.090 156.465 53.440 156.495 ;
        RECT 71.070 156.465 71.420 156.495 ;
        RECT 36.445 155.845 36.795 155.875 ;
        RECT 72.145 155.845 72.495 155.875 ;
        RECT 36.445 155.495 72.495 155.845 ;
        RECT 36.445 155.465 36.795 155.495 ;
        RECT 72.145 155.465 72.495 155.495 ;
        RECT 63.285 154.845 63.635 154.875 ;
        RECT 74.425 154.845 74.775 154.875 ;
        RECT 63.285 154.495 74.775 154.845 ;
        RECT 63.285 154.465 63.635 154.495 ;
        RECT 74.425 154.465 74.775 154.495 ;
        RECT 32.960 153.845 33.310 153.875 ;
        RECT 75.500 153.845 75.850 153.875 ;
        RECT 32.960 153.495 75.850 153.845 ;
        RECT 32.960 153.465 33.310 153.495 ;
        RECT 75.500 153.465 75.850 153.495 ;
        RECT 59.800 152.845 60.150 152.875 ;
        RECT 77.780 152.845 78.130 152.875 ;
        RECT 59.800 152.495 78.130 152.845 ;
        RECT 59.800 152.465 60.150 152.495 ;
        RECT 77.780 152.465 78.130 152.495 ;
        RECT 26.760 146.050 27.050 146.915 ;
        RECT 27.645 146.705 28.645 146.735 ;
        RECT 29.780 146.705 30.040 146.780 ;
        RECT 31.175 146.705 31.825 146.735 ;
        RECT 27.625 146.535 31.845 146.705 ;
        RECT 27.645 146.505 28.645 146.535 ;
        RECT 29.780 146.460 30.040 146.535 ;
        RECT 31.175 146.505 31.825 146.535 ;
        RECT 27.210 146.250 27.440 146.395 ;
        RECT 27.625 146.250 27.885 146.325 ;
        RECT 28.850 146.250 29.080 146.395 ;
        RECT 30.785 146.250 31.015 146.395 ;
        RECT 31.985 146.250 32.215 146.395 ;
        RECT 27.210 146.080 32.215 146.250 ;
        RECT 26.755 145.690 27.055 146.050 ;
        RECT 27.210 145.935 27.440 146.080 ;
        RECT 27.625 146.005 27.885 146.080 ;
        RECT 28.850 145.935 29.080 146.080 ;
        RECT 30.785 145.935 31.015 146.080 ;
        RECT 31.985 145.935 32.215 146.080 ;
        RECT 27.645 145.795 28.645 145.825 ;
        RECT 31.175 145.795 31.825 145.825 ;
        RECT 32.420 145.795 32.710 146.915 ;
        RECT 33.470 146.050 33.760 146.915 ;
        RECT 34.355 146.705 35.355 146.735 ;
        RECT 36.490 146.705 36.750 146.780 ;
        RECT 37.885 146.705 38.535 146.735 ;
        RECT 34.335 146.535 38.555 146.705 ;
        RECT 34.355 146.505 35.355 146.535 ;
        RECT 36.490 146.460 36.750 146.535 ;
        RECT 37.885 146.505 38.535 146.535 ;
        RECT 33.920 146.250 34.150 146.395 ;
        RECT 34.335 146.250 34.595 146.325 ;
        RECT 35.560 146.250 35.790 146.395 ;
        RECT 37.495 146.250 37.725 146.395 ;
        RECT 38.695 146.250 38.925 146.395 ;
        RECT 33.920 146.080 38.925 146.250 ;
        RECT 26.760 143.050 27.050 145.690 ;
        RECT 27.625 145.625 28.665 145.795 ;
        RECT 31.155 145.625 32.710 145.795 ;
        RECT 33.465 145.690 33.765 146.050 ;
        RECT 33.920 145.935 34.150 146.080 ;
        RECT 34.335 146.005 34.595 146.080 ;
        RECT 35.560 145.935 35.790 146.080 ;
        RECT 37.495 145.935 37.725 146.080 ;
        RECT 38.695 145.935 38.925 146.080 ;
        RECT 34.355 145.795 35.355 145.825 ;
        RECT 37.885 145.795 38.535 145.825 ;
        RECT 39.130 145.795 39.420 146.915 ;
        RECT 40.180 146.050 40.470 146.915 ;
        RECT 41.065 146.705 42.065 146.735 ;
        RECT 43.200 146.705 43.460 146.780 ;
        RECT 44.595 146.705 45.245 146.735 ;
        RECT 41.045 146.535 45.265 146.705 ;
        RECT 41.065 146.505 42.065 146.535 ;
        RECT 43.200 146.460 43.460 146.535 ;
        RECT 44.595 146.505 45.245 146.535 ;
        RECT 40.630 146.250 40.860 146.395 ;
        RECT 41.045 146.250 41.305 146.325 ;
        RECT 42.270 146.250 42.500 146.395 ;
        RECT 44.205 146.250 44.435 146.395 ;
        RECT 45.405 146.250 45.635 146.395 ;
        RECT 40.630 146.080 45.635 146.250 ;
        RECT 27.645 145.595 28.645 145.625 ;
        RECT 31.175 145.595 31.825 145.625 ;
        RECT 28.060 145.235 28.230 145.595 ;
        RECT 27.645 145.205 28.645 145.235 ;
        RECT 29.780 145.205 30.040 145.280 ;
        RECT 31.175 145.205 31.825 145.235 ;
        RECT 27.625 145.035 28.665 145.205 ;
        RECT 29.780 145.035 31.845 145.205 ;
        RECT 27.645 145.005 28.645 145.035 ;
        RECT 29.780 144.960 30.040 145.035 ;
        RECT 31.175 145.005 31.825 145.035 ;
        RECT 27.210 144.750 27.440 144.895 ;
        RECT 28.850 144.825 29.080 144.895 ;
        RECT 28.465 144.750 29.080 144.825 ;
        RECT 30.785 144.750 31.015 144.895 ;
        RECT 31.985 144.750 32.215 144.895 ;
        RECT 27.210 144.580 32.215 144.750 ;
        RECT 27.210 144.435 27.440 144.580 ;
        RECT 28.465 144.505 29.080 144.580 ;
        RECT 28.850 144.435 29.080 144.505 ;
        RECT 30.785 144.435 31.015 144.580 ;
        RECT 31.985 144.435 32.215 144.580 ;
        RECT 32.420 144.550 32.710 145.625 ;
        RECT 27.645 144.295 28.645 144.325 ;
        RECT 31.175 144.295 31.825 144.325 ;
        RECT 32.415 144.295 32.715 144.550 ;
        RECT 27.625 144.125 28.665 144.295 ;
        RECT 31.155 144.190 32.715 144.295 ;
        RECT 31.155 144.125 32.710 144.190 ;
        RECT 27.645 144.095 28.645 144.125 ;
        RECT 31.175 144.095 31.825 144.125 ;
        RECT 28.060 143.735 28.230 144.095 ;
        RECT 27.645 143.705 28.645 143.735 ;
        RECT 29.780 143.705 30.040 143.780 ;
        RECT 31.175 143.705 31.825 143.735 ;
        RECT 27.625 143.535 28.665 143.705 ;
        RECT 29.780 143.535 31.845 143.705 ;
        RECT 27.645 143.505 28.645 143.535 ;
        RECT 29.780 143.460 30.040 143.535 ;
        RECT 31.175 143.505 31.825 143.535 ;
        RECT 27.210 143.250 27.440 143.395 ;
        RECT 28.850 143.325 29.080 143.395 ;
        RECT 28.850 143.250 29.145 143.325 ;
        RECT 30.785 143.250 31.015 143.395 ;
        RECT 31.985 143.250 32.215 143.395 ;
        RECT 27.210 143.080 32.215 143.250 ;
        RECT 26.755 142.795 27.055 143.050 ;
        RECT 27.210 142.935 27.440 143.080 ;
        RECT 28.850 143.005 29.145 143.080 ;
        RECT 28.850 142.935 29.080 143.005 ;
        RECT 30.785 142.935 31.015 143.080 ;
        RECT 31.985 142.935 32.215 143.080 ;
        RECT 27.645 142.795 28.645 142.825 ;
        RECT 31.175 142.795 31.825 142.825 ;
        RECT 32.420 142.795 32.710 144.125 ;
        RECT 33.470 143.050 33.760 145.690 ;
        RECT 34.335 145.625 35.375 145.795 ;
        RECT 37.865 145.625 39.420 145.795 ;
        RECT 40.175 145.690 40.475 146.050 ;
        RECT 40.630 145.935 40.860 146.080 ;
        RECT 41.045 146.005 41.305 146.080 ;
        RECT 42.270 145.935 42.500 146.080 ;
        RECT 44.205 145.935 44.435 146.080 ;
        RECT 45.405 145.935 45.635 146.080 ;
        RECT 41.065 145.795 42.065 145.825 ;
        RECT 44.595 145.795 45.245 145.825 ;
        RECT 45.840 145.795 46.130 146.915 ;
        RECT 46.890 146.050 47.180 146.915 ;
        RECT 47.775 146.705 48.775 146.735 ;
        RECT 49.910 146.705 50.170 146.780 ;
        RECT 51.305 146.705 51.955 146.735 ;
        RECT 47.755 146.535 51.975 146.705 ;
        RECT 47.775 146.505 48.775 146.535 ;
        RECT 49.910 146.460 50.170 146.535 ;
        RECT 51.305 146.505 51.955 146.535 ;
        RECT 47.340 146.250 47.570 146.395 ;
        RECT 47.755 146.250 48.015 146.325 ;
        RECT 48.980 146.250 49.210 146.395 ;
        RECT 50.915 146.250 51.145 146.395 ;
        RECT 52.115 146.250 52.345 146.395 ;
        RECT 47.340 146.080 52.345 146.250 ;
        RECT 34.355 145.595 35.355 145.625 ;
        RECT 37.885 145.595 38.535 145.625 ;
        RECT 34.770 145.235 34.940 145.595 ;
        RECT 34.355 145.205 35.355 145.235 ;
        RECT 36.490 145.205 36.750 145.280 ;
        RECT 37.885 145.205 38.535 145.235 ;
        RECT 34.335 145.035 35.375 145.205 ;
        RECT 36.490 145.035 38.555 145.205 ;
        RECT 34.355 145.005 35.355 145.035 ;
        RECT 36.490 144.960 36.750 145.035 ;
        RECT 37.885 145.005 38.535 145.035 ;
        RECT 33.920 144.750 34.150 144.895 ;
        RECT 35.560 144.825 35.790 144.895 ;
        RECT 35.175 144.750 35.790 144.825 ;
        RECT 37.495 144.750 37.725 144.895 ;
        RECT 38.695 144.750 38.925 144.895 ;
        RECT 33.920 144.580 38.925 144.750 ;
        RECT 33.920 144.435 34.150 144.580 ;
        RECT 35.175 144.505 35.790 144.580 ;
        RECT 35.560 144.435 35.790 144.505 ;
        RECT 37.495 144.435 37.725 144.580 ;
        RECT 38.695 144.435 38.925 144.580 ;
        RECT 39.130 144.550 39.420 145.625 ;
        RECT 34.355 144.295 35.355 144.325 ;
        RECT 37.885 144.295 38.535 144.325 ;
        RECT 39.125 144.295 39.425 144.550 ;
        RECT 34.335 144.125 35.375 144.295 ;
        RECT 37.865 144.190 39.425 144.295 ;
        RECT 37.865 144.125 39.420 144.190 ;
        RECT 34.355 144.095 35.355 144.125 ;
        RECT 37.885 144.095 38.535 144.125 ;
        RECT 34.770 143.735 34.940 144.095 ;
        RECT 34.355 143.705 35.355 143.735 ;
        RECT 36.490 143.705 36.750 143.780 ;
        RECT 37.885 143.705 38.535 143.735 ;
        RECT 34.335 143.535 35.375 143.705 ;
        RECT 36.490 143.535 38.555 143.705 ;
        RECT 34.355 143.505 35.355 143.535 ;
        RECT 36.490 143.460 36.750 143.535 ;
        RECT 37.885 143.505 38.535 143.535 ;
        RECT 33.920 143.250 34.150 143.395 ;
        RECT 35.560 143.325 35.790 143.395 ;
        RECT 35.560 143.250 35.855 143.325 ;
        RECT 37.495 143.250 37.725 143.395 ;
        RECT 38.695 143.250 38.925 143.395 ;
        RECT 33.920 143.080 38.925 143.250 ;
        RECT 26.755 142.690 28.665 142.795 ;
        RECT 26.760 142.625 28.665 142.690 ;
        RECT 31.155 142.625 32.710 142.795 ;
        RECT 33.465 142.795 33.765 143.050 ;
        RECT 33.920 142.935 34.150 143.080 ;
        RECT 35.560 143.005 35.855 143.080 ;
        RECT 35.560 142.935 35.790 143.005 ;
        RECT 37.495 142.935 37.725 143.080 ;
        RECT 38.695 142.935 38.925 143.080 ;
        RECT 34.355 142.795 35.355 142.825 ;
        RECT 37.885 142.795 38.535 142.825 ;
        RECT 39.130 142.795 39.420 144.125 ;
        RECT 40.180 143.050 40.470 145.690 ;
        RECT 41.045 145.625 42.085 145.795 ;
        RECT 44.575 145.625 46.130 145.795 ;
        RECT 46.885 145.690 47.185 146.050 ;
        RECT 47.340 145.935 47.570 146.080 ;
        RECT 47.755 146.005 48.015 146.080 ;
        RECT 48.980 145.935 49.210 146.080 ;
        RECT 50.915 145.935 51.145 146.080 ;
        RECT 52.115 145.935 52.345 146.080 ;
        RECT 47.775 145.795 48.775 145.825 ;
        RECT 51.305 145.795 51.955 145.825 ;
        RECT 52.550 145.795 52.840 146.915 ;
        RECT 53.600 146.050 53.890 146.915 ;
        RECT 54.485 146.705 55.485 146.735 ;
        RECT 56.620 146.705 56.880 146.780 ;
        RECT 58.015 146.705 58.665 146.735 ;
        RECT 54.465 146.535 58.685 146.705 ;
        RECT 54.485 146.505 55.485 146.535 ;
        RECT 56.620 146.460 56.880 146.535 ;
        RECT 58.015 146.505 58.665 146.535 ;
        RECT 54.050 146.250 54.280 146.395 ;
        RECT 54.465 146.250 54.725 146.325 ;
        RECT 55.690 146.250 55.920 146.395 ;
        RECT 57.625 146.250 57.855 146.395 ;
        RECT 58.825 146.250 59.055 146.395 ;
        RECT 54.050 146.080 59.055 146.250 ;
        RECT 41.065 145.595 42.065 145.625 ;
        RECT 44.595 145.595 45.245 145.625 ;
        RECT 41.480 145.235 41.650 145.595 ;
        RECT 41.065 145.205 42.065 145.235 ;
        RECT 43.200 145.205 43.460 145.280 ;
        RECT 44.595 145.205 45.245 145.235 ;
        RECT 41.045 145.035 42.085 145.205 ;
        RECT 43.200 145.035 45.265 145.205 ;
        RECT 41.065 145.005 42.065 145.035 ;
        RECT 43.200 144.960 43.460 145.035 ;
        RECT 44.595 145.005 45.245 145.035 ;
        RECT 40.630 144.750 40.860 144.895 ;
        RECT 42.270 144.825 42.500 144.895 ;
        RECT 41.885 144.750 42.500 144.825 ;
        RECT 44.205 144.750 44.435 144.895 ;
        RECT 45.405 144.750 45.635 144.895 ;
        RECT 40.630 144.580 45.635 144.750 ;
        RECT 40.630 144.435 40.860 144.580 ;
        RECT 41.885 144.505 42.500 144.580 ;
        RECT 42.270 144.435 42.500 144.505 ;
        RECT 44.205 144.435 44.435 144.580 ;
        RECT 45.405 144.435 45.635 144.580 ;
        RECT 45.840 144.550 46.130 145.625 ;
        RECT 41.065 144.295 42.065 144.325 ;
        RECT 44.595 144.295 45.245 144.325 ;
        RECT 45.835 144.295 46.135 144.550 ;
        RECT 41.045 144.125 42.085 144.295 ;
        RECT 44.575 144.190 46.135 144.295 ;
        RECT 44.575 144.125 46.130 144.190 ;
        RECT 41.065 144.095 42.065 144.125 ;
        RECT 44.595 144.095 45.245 144.125 ;
        RECT 41.480 143.735 41.650 144.095 ;
        RECT 41.065 143.705 42.065 143.735 ;
        RECT 43.200 143.705 43.460 143.780 ;
        RECT 44.595 143.705 45.245 143.735 ;
        RECT 41.045 143.535 42.085 143.705 ;
        RECT 43.200 143.535 45.265 143.705 ;
        RECT 41.065 143.505 42.065 143.535 ;
        RECT 43.200 143.460 43.460 143.535 ;
        RECT 44.595 143.505 45.245 143.535 ;
        RECT 40.630 143.250 40.860 143.395 ;
        RECT 42.270 143.325 42.500 143.395 ;
        RECT 42.270 143.250 42.565 143.325 ;
        RECT 44.205 143.250 44.435 143.395 ;
        RECT 45.405 143.250 45.635 143.395 ;
        RECT 40.630 143.080 45.635 143.250 ;
        RECT 33.465 142.690 35.375 142.795 ;
        RECT 26.760 140.050 27.050 142.625 ;
        RECT 27.645 142.595 28.645 142.625 ;
        RECT 31.175 142.595 31.825 142.625 ;
        RECT 27.645 142.205 28.645 142.235 ;
        RECT 29.780 142.205 30.040 142.280 ;
        RECT 31.175 142.205 31.825 142.235 ;
        RECT 27.625 142.035 31.845 142.205 ;
        RECT 27.645 142.005 28.645 142.035 ;
        RECT 29.780 141.960 30.040 142.035 ;
        RECT 31.175 142.005 31.825 142.035 ;
        RECT 27.210 141.750 27.440 141.895 ;
        RECT 27.625 141.750 27.885 141.825 ;
        RECT 28.850 141.750 29.080 141.895 ;
        RECT 30.785 141.750 31.015 141.895 ;
        RECT 31.985 141.750 32.215 141.895 ;
        RECT 27.210 141.580 32.215 141.750 ;
        RECT 27.210 141.435 27.440 141.580 ;
        RECT 27.625 141.505 27.885 141.580 ;
        RECT 28.850 141.435 29.080 141.580 ;
        RECT 30.785 141.435 31.015 141.580 ;
        RECT 31.985 141.435 32.215 141.580 ;
        RECT 32.420 141.550 32.710 142.625 ;
        RECT 33.470 142.625 35.375 142.690 ;
        RECT 37.865 142.625 39.420 142.795 ;
        RECT 40.175 142.795 40.475 143.050 ;
        RECT 40.630 142.935 40.860 143.080 ;
        RECT 42.270 143.005 42.565 143.080 ;
        RECT 42.270 142.935 42.500 143.005 ;
        RECT 44.205 142.935 44.435 143.080 ;
        RECT 45.405 142.935 45.635 143.080 ;
        RECT 41.065 142.795 42.065 142.825 ;
        RECT 44.595 142.795 45.245 142.825 ;
        RECT 45.840 142.795 46.130 144.125 ;
        RECT 46.890 143.050 47.180 145.690 ;
        RECT 47.755 145.625 48.795 145.795 ;
        RECT 51.285 145.625 52.840 145.795 ;
        RECT 53.595 145.690 53.895 146.050 ;
        RECT 54.050 145.935 54.280 146.080 ;
        RECT 54.465 146.005 54.725 146.080 ;
        RECT 55.690 145.935 55.920 146.080 ;
        RECT 57.625 145.935 57.855 146.080 ;
        RECT 58.825 145.935 59.055 146.080 ;
        RECT 54.485 145.795 55.485 145.825 ;
        RECT 58.015 145.795 58.665 145.825 ;
        RECT 59.260 145.795 59.550 146.915 ;
        RECT 60.310 146.050 60.600 146.915 ;
        RECT 61.195 146.705 62.195 146.735 ;
        RECT 63.330 146.705 63.590 146.780 ;
        RECT 64.725 146.705 65.375 146.735 ;
        RECT 61.175 146.535 65.395 146.705 ;
        RECT 61.195 146.505 62.195 146.535 ;
        RECT 63.330 146.460 63.590 146.535 ;
        RECT 64.725 146.505 65.375 146.535 ;
        RECT 60.760 146.250 60.990 146.395 ;
        RECT 61.175 146.250 61.435 146.325 ;
        RECT 62.400 146.250 62.630 146.395 ;
        RECT 64.335 146.250 64.565 146.395 ;
        RECT 65.535 146.250 65.765 146.395 ;
        RECT 60.760 146.080 65.765 146.250 ;
        RECT 47.775 145.595 48.775 145.625 ;
        RECT 51.305 145.595 51.955 145.625 ;
        RECT 48.190 145.235 48.360 145.595 ;
        RECT 47.775 145.205 48.775 145.235 ;
        RECT 49.910 145.205 50.170 145.280 ;
        RECT 51.305 145.205 51.955 145.235 ;
        RECT 47.755 145.035 48.795 145.205 ;
        RECT 49.910 145.035 51.975 145.205 ;
        RECT 47.775 145.005 48.775 145.035 ;
        RECT 49.910 144.960 50.170 145.035 ;
        RECT 51.305 145.005 51.955 145.035 ;
        RECT 47.340 144.750 47.570 144.895 ;
        RECT 48.980 144.825 49.210 144.895 ;
        RECT 48.595 144.750 49.210 144.825 ;
        RECT 50.915 144.750 51.145 144.895 ;
        RECT 52.115 144.750 52.345 144.895 ;
        RECT 47.340 144.580 52.345 144.750 ;
        RECT 47.340 144.435 47.570 144.580 ;
        RECT 48.595 144.505 49.210 144.580 ;
        RECT 48.980 144.435 49.210 144.505 ;
        RECT 50.915 144.435 51.145 144.580 ;
        RECT 52.115 144.435 52.345 144.580 ;
        RECT 52.550 144.550 52.840 145.625 ;
        RECT 47.775 144.295 48.775 144.325 ;
        RECT 51.305 144.295 51.955 144.325 ;
        RECT 52.545 144.295 52.845 144.550 ;
        RECT 47.755 144.125 48.795 144.295 ;
        RECT 51.285 144.190 52.845 144.295 ;
        RECT 51.285 144.125 52.840 144.190 ;
        RECT 47.775 144.095 48.775 144.125 ;
        RECT 51.305 144.095 51.955 144.125 ;
        RECT 48.190 143.735 48.360 144.095 ;
        RECT 47.775 143.705 48.775 143.735 ;
        RECT 49.910 143.705 50.170 143.780 ;
        RECT 51.305 143.705 51.955 143.735 ;
        RECT 47.755 143.535 48.795 143.705 ;
        RECT 49.910 143.535 51.975 143.705 ;
        RECT 47.775 143.505 48.775 143.535 ;
        RECT 49.910 143.460 50.170 143.535 ;
        RECT 51.305 143.505 51.955 143.535 ;
        RECT 47.340 143.250 47.570 143.395 ;
        RECT 48.980 143.325 49.210 143.395 ;
        RECT 48.980 143.250 49.275 143.325 ;
        RECT 50.915 143.250 51.145 143.395 ;
        RECT 52.115 143.250 52.345 143.395 ;
        RECT 47.340 143.080 52.345 143.250 ;
        RECT 40.175 142.690 42.085 142.795 ;
        RECT 27.645 141.295 28.645 141.325 ;
        RECT 31.175 141.295 31.825 141.325 ;
        RECT 32.415 141.295 32.715 141.550 ;
        RECT 27.625 141.125 28.665 141.295 ;
        RECT 31.155 141.190 32.715 141.295 ;
        RECT 31.155 141.125 32.710 141.190 ;
        RECT 27.645 141.095 28.645 141.125 ;
        RECT 31.175 141.095 31.825 141.125 ;
        RECT 28.060 140.735 28.230 141.095 ;
        RECT 27.645 140.705 28.645 140.735 ;
        RECT 29.780 140.705 30.040 140.780 ;
        RECT 31.175 140.705 31.825 140.735 ;
        RECT 27.625 140.535 28.665 140.705 ;
        RECT 29.780 140.535 31.845 140.705 ;
        RECT 27.645 140.505 28.645 140.535 ;
        RECT 29.780 140.460 30.040 140.535 ;
        RECT 31.175 140.505 31.825 140.535 ;
        RECT 27.210 140.250 27.440 140.395 ;
        RECT 28.045 140.250 28.305 140.325 ;
        RECT 28.850 140.250 29.080 140.395 ;
        RECT 30.785 140.250 31.015 140.395 ;
        RECT 31.985 140.250 32.215 140.395 ;
        RECT 27.210 140.080 32.215 140.250 ;
        RECT 26.755 139.690 27.055 140.050 ;
        RECT 27.210 139.935 27.440 140.080 ;
        RECT 28.045 140.005 28.305 140.080 ;
        RECT 28.850 139.935 29.080 140.080 ;
        RECT 30.785 139.935 31.015 140.080 ;
        RECT 31.985 139.935 32.215 140.080 ;
        RECT 27.645 139.795 28.645 139.825 ;
        RECT 31.175 139.795 31.825 139.825 ;
        RECT 32.420 139.795 32.710 141.125 ;
        RECT 33.470 140.050 33.760 142.625 ;
        RECT 34.355 142.595 35.355 142.625 ;
        RECT 37.885 142.595 38.535 142.625 ;
        RECT 34.355 142.205 35.355 142.235 ;
        RECT 36.490 142.205 36.750 142.280 ;
        RECT 37.885 142.205 38.535 142.235 ;
        RECT 34.335 142.035 38.555 142.205 ;
        RECT 34.355 142.005 35.355 142.035 ;
        RECT 36.490 141.960 36.750 142.035 ;
        RECT 37.885 142.005 38.535 142.035 ;
        RECT 33.920 141.750 34.150 141.895 ;
        RECT 34.335 141.750 34.595 141.825 ;
        RECT 35.560 141.750 35.790 141.895 ;
        RECT 37.495 141.750 37.725 141.895 ;
        RECT 38.695 141.750 38.925 141.895 ;
        RECT 33.920 141.580 38.925 141.750 ;
        RECT 33.920 141.435 34.150 141.580 ;
        RECT 34.335 141.505 34.595 141.580 ;
        RECT 35.560 141.435 35.790 141.580 ;
        RECT 37.495 141.435 37.725 141.580 ;
        RECT 38.695 141.435 38.925 141.580 ;
        RECT 39.130 141.550 39.420 142.625 ;
        RECT 40.180 142.625 42.085 142.690 ;
        RECT 44.575 142.625 46.130 142.795 ;
        RECT 46.885 142.795 47.185 143.050 ;
        RECT 47.340 142.935 47.570 143.080 ;
        RECT 48.980 143.005 49.275 143.080 ;
        RECT 48.980 142.935 49.210 143.005 ;
        RECT 50.915 142.935 51.145 143.080 ;
        RECT 52.115 142.935 52.345 143.080 ;
        RECT 47.775 142.795 48.775 142.825 ;
        RECT 51.305 142.795 51.955 142.825 ;
        RECT 52.550 142.795 52.840 144.125 ;
        RECT 53.600 143.050 53.890 145.690 ;
        RECT 54.465 145.625 55.505 145.795 ;
        RECT 57.995 145.625 59.550 145.795 ;
        RECT 60.305 145.690 60.605 146.050 ;
        RECT 60.760 145.935 60.990 146.080 ;
        RECT 61.175 146.005 61.435 146.080 ;
        RECT 62.400 145.935 62.630 146.080 ;
        RECT 64.335 145.935 64.565 146.080 ;
        RECT 65.535 145.935 65.765 146.080 ;
        RECT 61.195 145.795 62.195 145.825 ;
        RECT 64.725 145.795 65.375 145.825 ;
        RECT 65.970 145.795 66.260 146.915 ;
        RECT 67.020 146.050 67.310 146.915 ;
        RECT 67.905 146.705 68.905 146.735 ;
        RECT 70.040 146.705 70.300 146.780 ;
        RECT 71.435 146.705 72.085 146.735 ;
        RECT 67.885 146.535 72.105 146.705 ;
        RECT 67.905 146.505 68.905 146.535 ;
        RECT 70.040 146.460 70.300 146.535 ;
        RECT 71.435 146.505 72.085 146.535 ;
        RECT 67.470 146.250 67.700 146.395 ;
        RECT 67.885 146.250 68.145 146.325 ;
        RECT 69.110 146.250 69.340 146.395 ;
        RECT 71.045 146.250 71.275 146.395 ;
        RECT 72.245 146.250 72.475 146.395 ;
        RECT 67.470 146.080 72.475 146.250 ;
        RECT 54.485 145.595 55.485 145.625 ;
        RECT 58.015 145.595 58.665 145.625 ;
        RECT 54.900 145.235 55.070 145.595 ;
        RECT 54.485 145.205 55.485 145.235 ;
        RECT 56.620 145.205 56.880 145.280 ;
        RECT 58.015 145.205 58.665 145.235 ;
        RECT 54.465 145.035 55.505 145.205 ;
        RECT 56.620 145.035 58.685 145.205 ;
        RECT 54.485 145.005 55.485 145.035 ;
        RECT 56.620 144.960 56.880 145.035 ;
        RECT 58.015 145.005 58.665 145.035 ;
        RECT 54.050 144.750 54.280 144.895 ;
        RECT 55.690 144.825 55.920 144.895 ;
        RECT 55.305 144.750 55.920 144.825 ;
        RECT 57.625 144.750 57.855 144.895 ;
        RECT 58.825 144.750 59.055 144.895 ;
        RECT 54.050 144.580 59.055 144.750 ;
        RECT 54.050 144.435 54.280 144.580 ;
        RECT 55.305 144.505 55.920 144.580 ;
        RECT 55.690 144.435 55.920 144.505 ;
        RECT 57.625 144.435 57.855 144.580 ;
        RECT 58.825 144.435 59.055 144.580 ;
        RECT 59.260 144.550 59.550 145.625 ;
        RECT 54.485 144.295 55.485 144.325 ;
        RECT 58.015 144.295 58.665 144.325 ;
        RECT 59.255 144.295 59.555 144.550 ;
        RECT 54.465 144.125 55.505 144.295 ;
        RECT 57.995 144.190 59.555 144.295 ;
        RECT 57.995 144.125 59.550 144.190 ;
        RECT 54.485 144.095 55.485 144.125 ;
        RECT 58.015 144.095 58.665 144.125 ;
        RECT 54.900 143.735 55.070 144.095 ;
        RECT 54.485 143.705 55.485 143.735 ;
        RECT 56.620 143.705 56.880 143.780 ;
        RECT 58.015 143.705 58.665 143.735 ;
        RECT 54.465 143.535 55.505 143.705 ;
        RECT 56.620 143.535 58.685 143.705 ;
        RECT 54.485 143.505 55.485 143.535 ;
        RECT 56.620 143.460 56.880 143.535 ;
        RECT 58.015 143.505 58.665 143.535 ;
        RECT 54.050 143.250 54.280 143.395 ;
        RECT 55.690 143.325 55.920 143.395 ;
        RECT 55.690 143.250 55.985 143.325 ;
        RECT 57.625 143.250 57.855 143.395 ;
        RECT 58.825 143.250 59.055 143.395 ;
        RECT 54.050 143.080 59.055 143.250 ;
        RECT 46.885 142.690 48.795 142.795 ;
        RECT 34.355 141.295 35.355 141.325 ;
        RECT 37.885 141.295 38.535 141.325 ;
        RECT 39.125 141.295 39.425 141.550 ;
        RECT 34.335 141.125 35.375 141.295 ;
        RECT 37.865 141.190 39.425 141.295 ;
        RECT 37.865 141.125 39.420 141.190 ;
        RECT 34.355 141.095 35.355 141.125 ;
        RECT 37.885 141.095 38.535 141.125 ;
        RECT 34.770 140.735 34.940 141.095 ;
        RECT 34.355 140.705 35.355 140.735 ;
        RECT 36.490 140.705 36.750 140.780 ;
        RECT 37.885 140.705 38.535 140.735 ;
        RECT 34.335 140.535 35.375 140.705 ;
        RECT 36.490 140.535 38.555 140.705 ;
        RECT 34.355 140.505 35.355 140.535 ;
        RECT 36.490 140.460 36.750 140.535 ;
        RECT 37.885 140.505 38.535 140.535 ;
        RECT 33.920 140.250 34.150 140.395 ;
        RECT 34.755 140.250 35.015 140.325 ;
        RECT 35.560 140.250 35.790 140.395 ;
        RECT 37.495 140.250 37.725 140.395 ;
        RECT 38.695 140.250 38.925 140.395 ;
        RECT 33.920 140.080 38.925 140.250 ;
        RECT 26.760 138.295 27.050 139.690 ;
        RECT 27.625 139.625 28.665 139.795 ;
        RECT 31.155 139.625 32.710 139.795 ;
        RECT 33.465 139.690 33.765 140.050 ;
        RECT 33.920 139.935 34.150 140.080 ;
        RECT 34.755 140.005 35.015 140.080 ;
        RECT 35.560 139.935 35.790 140.080 ;
        RECT 37.495 139.935 37.725 140.080 ;
        RECT 38.695 139.935 38.925 140.080 ;
        RECT 34.355 139.795 35.355 139.825 ;
        RECT 37.885 139.795 38.535 139.825 ;
        RECT 39.130 139.795 39.420 141.125 ;
        RECT 40.180 140.050 40.470 142.625 ;
        RECT 41.065 142.595 42.065 142.625 ;
        RECT 44.595 142.595 45.245 142.625 ;
        RECT 41.065 142.205 42.065 142.235 ;
        RECT 43.200 142.205 43.460 142.280 ;
        RECT 44.595 142.205 45.245 142.235 ;
        RECT 41.045 142.035 45.265 142.205 ;
        RECT 41.065 142.005 42.065 142.035 ;
        RECT 43.200 141.960 43.460 142.035 ;
        RECT 44.595 142.005 45.245 142.035 ;
        RECT 40.630 141.750 40.860 141.895 ;
        RECT 41.045 141.750 41.305 141.825 ;
        RECT 42.270 141.750 42.500 141.895 ;
        RECT 44.205 141.750 44.435 141.895 ;
        RECT 45.405 141.750 45.635 141.895 ;
        RECT 40.630 141.580 45.635 141.750 ;
        RECT 40.630 141.435 40.860 141.580 ;
        RECT 41.045 141.505 41.305 141.580 ;
        RECT 42.270 141.435 42.500 141.580 ;
        RECT 44.205 141.435 44.435 141.580 ;
        RECT 45.405 141.435 45.635 141.580 ;
        RECT 45.840 141.550 46.130 142.625 ;
        RECT 46.890 142.625 48.795 142.690 ;
        RECT 51.285 142.625 52.840 142.795 ;
        RECT 53.595 142.795 53.895 143.050 ;
        RECT 54.050 142.935 54.280 143.080 ;
        RECT 55.690 143.005 55.985 143.080 ;
        RECT 55.690 142.935 55.920 143.005 ;
        RECT 57.625 142.935 57.855 143.080 ;
        RECT 58.825 142.935 59.055 143.080 ;
        RECT 54.485 142.795 55.485 142.825 ;
        RECT 58.015 142.795 58.665 142.825 ;
        RECT 59.260 142.795 59.550 144.125 ;
        RECT 60.310 143.050 60.600 145.690 ;
        RECT 61.175 145.625 62.215 145.795 ;
        RECT 64.705 145.625 66.260 145.795 ;
        RECT 67.015 145.690 67.315 146.050 ;
        RECT 67.470 145.935 67.700 146.080 ;
        RECT 67.885 146.005 68.145 146.080 ;
        RECT 69.110 145.935 69.340 146.080 ;
        RECT 71.045 145.935 71.275 146.080 ;
        RECT 72.245 145.935 72.475 146.080 ;
        RECT 67.905 145.795 68.905 145.825 ;
        RECT 71.435 145.795 72.085 145.825 ;
        RECT 72.680 145.795 72.970 146.915 ;
        RECT 73.730 146.050 74.020 146.915 ;
        RECT 74.615 146.705 75.615 146.735 ;
        RECT 76.750 146.705 77.010 146.780 ;
        RECT 78.145 146.705 78.795 146.735 ;
        RECT 74.595 146.535 78.815 146.705 ;
        RECT 74.615 146.505 75.615 146.535 ;
        RECT 76.750 146.460 77.010 146.535 ;
        RECT 78.145 146.505 78.795 146.535 ;
        RECT 74.180 146.250 74.410 146.395 ;
        RECT 74.595 146.250 74.855 146.325 ;
        RECT 75.820 146.250 76.050 146.395 ;
        RECT 77.755 146.250 77.985 146.395 ;
        RECT 78.955 146.250 79.185 146.395 ;
        RECT 74.180 146.080 79.185 146.250 ;
        RECT 61.195 145.595 62.195 145.625 ;
        RECT 64.725 145.595 65.375 145.625 ;
        RECT 61.610 145.235 61.780 145.595 ;
        RECT 61.195 145.205 62.195 145.235 ;
        RECT 63.330 145.205 63.590 145.280 ;
        RECT 64.725 145.205 65.375 145.235 ;
        RECT 61.175 145.035 62.215 145.205 ;
        RECT 63.330 145.035 65.395 145.205 ;
        RECT 61.195 145.005 62.195 145.035 ;
        RECT 63.330 144.960 63.590 145.035 ;
        RECT 64.725 145.005 65.375 145.035 ;
        RECT 60.760 144.750 60.990 144.895 ;
        RECT 62.400 144.825 62.630 144.895 ;
        RECT 62.015 144.750 62.630 144.825 ;
        RECT 64.335 144.750 64.565 144.895 ;
        RECT 65.535 144.750 65.765 144.895 ;
        RECT 60.760 144.580 65.765 144.750 ;
        RECT 60.760 144.435 60.990 144.580 ;
        RECT 62.015 144.505 62.630 144.580 ;
        RECT 62.400 144.435 62.630 144.505 ;
        RECT 64.335 144.435 64.565 144.580 ;
        RECT 65.535 144.435 65.765 144.580 ;
        RECT 65.970 144.550 66.260 145.625 ;
        RECT 61.195 144.295 62.195 144.325 ;
        RECT 64.725 144.295 65.375 144.325 ;
        RECT 65.965 144.295 66.265 144.550 ;
        RECT 61.175 144.125 62.215 144.295 ;
        RECT 64.705 144.190 66.265 144.295 ;
        RECT 64.705 144.125 66.260 144.190 ;
        RECT 61.195 144.095 62.195 144.125 ;
        RECT 64.725 144.095 65.375 144.125 ;
        RECT 61.610 143.735 61.780 144.095 ;
        RECT 61.195 143.705 62.195 143.735 ;
        RECT 63.330 143.705 63.590 143.780 ;
        RECT 64.725 143.705 65.375 143.735 ;
        RECT 61.175 143.535 62.215 143.705 ;
        RECT 63.330 143.535 65.395 143.705 ;
        RECT 61.195 143.505 62.195 143.535 ;
        RECT 63.330 143.460 63.590 143.535 ;
        RECT 64.725 143.505 65.375 143.535 ;
        RECT 60.760 143.250 60.990 143.395 ;
        RECT 62.400 143.325 62.630 143.395 ;
        RECT 62.400 143.250 62.695 143.325 ;
        RECT 64.335 143.250 64.565 143.395 ;
        RECT 65.535 143.250 65.765 143.395 ;
        RECT 60.760 143.080 65.765 143.250 ;
        RECT 53.595 142.690 55.505 142.795 ;
        RECT 41.065 141.295 42.065 141.325 ;
        RECT 44.595 141.295 45.245 141.325 ;
        RECT 45.835 141.295 46.135 141.550 ;
        RECT 41.045 141.125 42.085 141.295 ;
        RECT 44.575 141.190 46.135 141.295 ;
        RECT 44.575 141.125 46.130 141.190 ;
        RECT 41.065 141.095 42.065 141.125 ;
        RECT 44.595 141.095 45.245 141.125 ;
        RECT 41.480 140.735 41.650 141.095 ;
        RECT 41.065 140.705 42.065 140.735 ;
        RECT 43.200 140.705 43.460 140.780 ;
        RECT 44.595 140.705 45.245 140.735 ;
        RECT 41.045 140.535 42.085 140.705 ;
        RECT 43.200 140.535 45.265 140.705 ;
        RECT 41.065 140.505 42.065 140.535 ;
        RECT 43.200 140.460 43.460 140.535 ;
        RECT 44.595 140.505 45.245 140.535 ;
        RECT 40.630 140.250 40.860 140.395 ;
        RECT 41.465 140.250 41.725 140.325 ;
        RECT 42.270 140.250 42.500 140.395 ;
        RECT 44.205 140.250 44.435 140.395 ;
        RECT 45.405 140.250 45.635 140.395 ;
        RECT 40.630 140.080 45.635 140.250 ;
        RECT 27.645 139.595 28.645 139.625 ;
        RECT 31.175 139.595 31.825 139.625 ;
        RECT 28.060 139.235 28.230 139.595 ;
        RECT 27.645 139.205 28.645 139.235 ;
        RECT 29.780 139.205 30.040 139.280 ;
        RECT 31.175 139.205 31.825 139.235 ;
        RECT 27.625 139.035 28.665 139.205 ;
        RECT 29.780 139.035 31.845 139.205 ;
        RECT 27.645 139.005 28.645 139.035 ;
        RECT 29.780 138.960 30.040 139.035 ;
        RECT 31.175 139.005 31.825 139.035 ;
        RECT 27.210 138.750 27.440 138.895 ;
        RECT 28.850 138.825 29.080 138.895 ;
        RECT 28.850 138.750 29.145 138.825 ;
        RECT 30.785 138.750 31.015 138.895 ;
        RECT 31.985 138.750 32.215 138.895 ;
        RECT 27.210 138.580 32.215 138.750 ;
        RECT 27.210 138.435 27.440 138.580 ;
        RECT 28.850 138.505 29.145 138.580 ;
        RECT 28.850 138.435 29.080 138.505 ;
        RECT 30.785 138.435 31.015 138.580 ;
        RECT 31.985 138.435 32.215 138.580 ;
        RECT 32.420 138.550 32.710 139.625 ;
        RECT 27.645 138.295 28.645 138.325 ;
        RECT 31.175 138.295 31.825 138.325 ;
        RECT 32.415 138.295 32.715 138.550 ;
        RECT 26.760 138.125 28.665 138.295 ;
        RECT 31.155 138.190 32.715 138.295 ;
        RECT 33.470 138.295 33.760 139.690 ;
        RECT 34.335 139.625 35.375 139.795 ;
        RECT 37.865 139.625 39.420 139.795 ;
        RECT 40.175 139.690 40.475 140.050 ;
        RECT 40.630 139.935 40.860 140.080 ;
        RECT 41.465 140.005 41.725 140.080 ;
        RECT 42.270 139.935 42.500 140.080 ;
        RECT 44.205 139.935 44.435 140.080 ;
        RECT 45.405 139.935 45.635 140.080 ;
        RECT 41.065 139.795 42.065 139.825 ;
        RECT 44.595 139.795 45.245 139.825 ;
        RECT 45.840 139.795 46.130 141.125 ;
        RECT 46.890 140.050 47.180 142.625 ;
        RECT 47.775 142.595 48.775 142.625 ;
        RECT 51.305 142.595 51.955 142.625 ;
        RECT 47.775 142.205 48.775 142.235 ;
        RECT 49.910 142.205 50.170 142.280 ;
        RECT 51.305 142.205 51.955 142.235 ;
        RECT 47.755 142.035 51.975 142.205 ;
        RECT 47.775 142.005 48.775 142.035 ;
        RECT 49.910 141.960 50.170 142.035 ;
        RECT 51.305 142.005 51.955 142.035 ;
        RECT 47.340 141.750 47.570 141.895 ;
        RECT 47.755 141.750 48.015 141.825 ;
        RECT 48.980 141.750 49.210 141.895 ;
        RECT 50.915 141.750 51.145 141.895 ;
        RECT 52.115 141.750 52.345 141.895 ;
        RECT 47.340 141.580 52.345 141.750 ;
        RECT 47.340 141.435 47.570 141.580 ;
        RECT 47.755 141.505 48.015 141.580 ;
        RECT 48.980 141.435 49.210 141.580 ;
        RECT 50.915 141.435 51.145 141.580 ;
        RECT 52.115 141.435 52.345 141.580 ;
        RECT 52.550 141.550 52.840 142.625 ;
        RECT 53.600 142.625 55.505 142.690 ;
        RECT 57.995 142.625 59.550 142.795 ;
        RECT 60.305 142.795 60.605 143.050 ;
        RECT 60.760 142.935 60.990 143.080 ;
        RECT 62.400 143.005 62.695 143.080 ;
        RECT 62.400 142.935 62.630 143.005 ;
        RECT 64.335 142.935 64.565 143.080 ;
        RECT 65.535 142.935 65.765 143.080 ;
        RECT 61.195 142.795 62.195 142.825 ;
        RECT 64.725 142.795 65.375 142.825 ;
        RECT 65.970 142.795 66.260 144.125 ;
        RECT 67.020 143.050 67.310 145.690 ;
        RECT 67.885 145.625 68.925 145.795 ;
        RECT 71.415 145.625 72.970 145.795 ;
        RECT 73.725 145.690 74.025 146.050 ;
        RECT 74.180 145.935 74.410 146.080 ;
        RECT 74.595 146.005 74.855 146.080 ;
        RECT 75.820 145.935 76.050 146.080 ;
        RECT 77.755 145.935 77.985 146.080 ;
        RECT 78.955 145.935 79.185 146.080 ;
        RECT 74.615 145.795 75.615 145.825 ;
        RECT 78.145 145.795 78.795 145.825 ;
        RECT 79.390 145.795 79.680 146.915 ;
        RECT 80.440 146.050 80.730 146.915 ;
        RECT 81.325 146.705 82.325 146.735 ;
        RECT 83.460 146.705 83.720 146.780 ;
        RECT 84.855 146.705 85.505 146.735 ;
        RECT 81.305 146.535 85.525 146.705 ;
        RECT 81.325 146.505 82.325 146.535 ;
        RECT 83.460 146.460 83.720 146.535 ;
        RECT 84.855 146.505 85.505 146.535 ;
        RECT 80.890 146.250 81.120 146.395 ;
        RECT 81.305 146.250 81.565 146.325 ;
        RECT 82.530 146.250 82.760 146.395 ;
        RECT 84.465 146.250 84.695 146.395 ;
        RECT 85.665 146.250 85.895 146.395 ;
        RECT 80.890 146.080 85.895 146.250 ;
        RECT 67.905 145.595 68.905 145.625 ;
        RECT 71.435 145.595 72.085 145.625 ;
        RECT 68.320 145.235 68.490 145.595 ;
        RECT 67.905 145.205 68.905 145.235 ;
        RECT 70.040 145.205 70.300 145.280 ;
        RECT 71.435 145.205 72.085 145.235 ;
        RECT 67.885 145.035 68.925 145.205 ;
        RECT 70.040 145.035 72.105 145.205 ;
        RECT 67.905 145.005 68.905 145.035 ;
        RECT 70.040 144.960 70.300 145.035 ;
        RECT 71.435 145.005 72.085 145.035 ;
        RECT 67.470 144.750 67.700 144.895 ;
        RECT 69.110 144.825 69.340 144.895 ;
        RECT 68.725 144.750 69.340 144.825 ;
        RECT 71.045 144.750 71.275 144.895 ;
        RECT 72.245 144.750 72.475 144.895 ;
        RECT 67.470 144.580 72.475 144.750 ;
        RECT 67.470 144.435 67.700 144.580 ;
        RECT 68.725 144.505 69.340 144.580 ;
        RECT 69.110 144.435 69.340 144.505 ;
        RECT 71.045 144.435 71.275 144.580 ;
        RECT 72.245 144.435 72.475 144.580 ;
        RECT 72.680 144.550 72.970 145.625 ;
        RECT 67.905 144.295 68.905 144.325 ;
        RECT 71.435 144.295 72.085 144.325 ;
        RECT 72.675 144.295 72.975 144.550 ;
        RECT 67.885 144.125 68.925 144.295 ;
        RECT 71.415 144.190 72.975 144.295 ;
        RECT 71.415 144.125 72.970 144.190 ;
        RECT 67.905 144.095 68.905 144.125 ;
        RECT 71.435 144.095 72.085 144.125 ;
        RECT 68.320 143.735 68.490 144.095 ;
        RECT 67.905 143.705 68.905 143.735 ;
        RECT 70.040 143.705 70.300 143.780 ;
        RECT 71.435 143.705 72.085 143.735 ;
        RECT 67.885 143.535 68.925 143.705 ;
        RECT 70.040 143.535 72.105 143.705 ;
        RECT 67.905 143.505 68.905 143.535 ;
        RECT 70.040 143.460 70.300 143.535 ;
        RECT 71.435 143.505 72.085 143.535 ;
        RECT 67.470 143.250 67.700 143.395 ;
        RECT 69.110 143.325 69.340 143.395 ;
        RECT 69.110 143.250 69.405 143.325 ;
        RECT 71.045 143.250 71.275 143.395 ;
        RECT 72.245 143.250 72.475 143.395 ;
        RECT 67.470 143.080 72.475 143.250 ;
        RECT 60.305 142.690 62.215 142.795 ;
        RECT 47.775 141.295 48.775 141.325 ;
        RECT 51.305 141.295 51.955 141.325 ;
        RECT 52.545 141.295 52.845 141.550 ;
        RECT 47.755 141.125 48.795 141.295 ;
        RECT 51.285 141.190 52.845 141.295 ;
        RECT 51.285 141.125 52.840 141.190 ;
        RECT 47.775 141.095 48.775 141.125 ;
        RECT 51.305 141.095 51.955 141.125 ;
        RECT 48.190 140.735 48.360 141.095 ;
        RECT 47.775 140.705 48.775 140.735 ;
        RECT 49.910 140.705 50.170 140.780 ;
        RECT 51.305 140.705 51.955 140.735 ;
        RECT 47.755 140.535 48.795 140.705 ;
        RECT 49.910 140.535 51.975 140.705 ;
        RECT 47.775 140.505 48.775 140.535 ;
        RECT 49.910 140.460 50.170 140.535 ;
        RECT 51.305 140.505 51.955 140.535 ;
        RECT 47.340 140.250 47.570 140.395 ;
        RECT 48.175 140.250 48.435 140.325 ;
        RECT 48.980 140.250 49.210 140.395 ;
        RECT 50.915 140.250 51.145 140.395 ;
        RECT 52.115 140.250 52.345 140.395 ;
        RECT 47.340 140.080 52.345 140.250 ;
        RECT 34.355 139.595 35.355 139.625 ;
        RECT 37.885 139.595 38.535 139.625 ;
        RECT 34.770 139.235 34.940 139.595 ;
        RECT 34.355 139.205 35.355 139.235 ;
        RECT 36.490 139.205 36.750 139.280 ;
        RECT 37.885 139.205 38.535 139.235 ;
        RECT 34.335 139.035 35.375 139.205 ;
        RECT 36.490 139.035 38.555 139.205 ;
        RECT 34.355 139.005 35.355 139.035 ;
        RECT 36.490 138.960 36.750 139.035 ;
        RECT 37.885 139.005 38.535 139.035 ;
        RECT 33.920 138.750 34.150 138.895 ;
        RECT 35.560 138.825 35.790 138.895 ;
        RECT 35.560 138.750 35.855 138.825 ;
        RECT 37.495 138.750 37.725 138.895 ;
        RECT 38.695 138.750 38.925 138.895 ;
        RECT 33.920 138.580 38.925 138.750 ;
        RECT 33.920 138.435 34.150 138.580 ;
        RECT 35.560 138.505 35.855 138.580 ;
        RECT 35.560 138.435 35.790 138.505 ;
        RECT 37.495 138.435 37.725 138.580 ;
        RECT 38.695 138.435 38.925 138.580 ;
        RECT 39.130 138.550 39.420 139.625 ;
        RECT 34.355 138.295 35.355 138.325 ;
        RECT 37.885 138.295 38.535 138.325 ;
        RECT 39.125 138.295 39.425 138.550 ;
        RECT 31.155 138.125 32.710 138.190 ;
        RECT 26.760 137.050 27.050 138.125 ;
        RECT 27.645 138.095 28.645 138.125 ;
        RECT 31.175 138.095 31.825 138.125 ;
        RECT 31.585 137.735 31.845 137.780 ;
        RECT 27.645 137.705 28.645 137.735 ;
        RECT 31.175 137.705 31.845 137.735 ;
        RECT 27.625 137.535 31.845 137.705 ;
        RECT 27.645 137.505 28.645 137.535 ;
        RECT 31.175 137.505 31.845 137.535 ;
        RECT 31.585 137.460 31.845 137.505 ;
        RECT 27.210 137.250 27.440 137.395 ;
        RECT 28.850 137.250 29.080 137.395 ;
        RECT 29.780 137.250 30.040 137.325 ;
        RECT 30.785 137.250 31.015 137.395 ;
        RECT 31.985 137.250 32.215 137.395 ;
        RECT 27.210 137.080 32.215 137.250 ;
        RECT 26.755 136.795 27.055 137.050 ;
        RECT 27.210 136.935 27.440 137.080 ;
        RECT 28.850 136.935 29.080 137.080 ;
        RECT 29.780 137.005 30.040 137.080 ;
        RECT 30.785 136.935 31.015 137.080 ;
        RECT 31.985 136.935 32.215 137.080 ;
        RECT 27.645 136.795 28.645 136.825 ;
        RECT 31.175 136.795 31.825 136.825 ;
        RECT 32.420 136.795 32.710 138.125 ;
        RECT 33.470 138.125 35.375 138.295 ;
        RECT 37.865 138.190 39.425 138.295 ;
        RECT 40.180 138.295 40.470 139.690 ;
        RECT 41.045 139.625 42.085 139.795 ;
        RECT 44.575 139.625 46.130 139.795 ;
        RECT 46.885 139.690 47.185 140.050 ;
        RECT 47.340 139.935 47.570 140.080 ;
        RECT 48.175 140.005 48.435 140.080 ;
        RECT 48.980 139.935 49.210 140.080 ;
        RECT 50.915 139.935 51.145 140.080 ;
        RECT 52.115 139.935 52.345 140.080 ;
        RECT 47.775 139.795 48.775 139.825 ;
        RECT 51.305 139.795 51.955 139.825 ;
        RECT 52.550 139.795 52.840 141.125 ;
        RECT 53.600 140.050 53.890 142.625 ;
        RECT 54.485 142.595 55.485 142.625 ;
        RECT 58.015 142.595 58.665 142.625 ;
        RECT 54.485 142.205 55.485 142.235 ;
        RECT 56.620 142.205 56.880 142.280 ;
        RECT 58.015 142.205 58.665 142.235 ;
        RECT 54.465 142.035 58.685 142.205 ;
        RECT 54.485 142.005 55.485 142.035 ;
        RECT 56.620 141.960 56.880 142.035 ;
        RECT 58.015 142.005 58.665 142.035 ;
        RECT 54.050 141.750 54.280 141.895 ;
        RECT 54.465 141.750 54.725 141.825 ;
        RECT 55.690 141.750 55.920 141.895 ;
        RECT 57.625 141.750 57.855 141.895 ;
        RECT 58.825 141.750 59.055 141.895 ;
        RECT 54.050 141.580 59.055 141.750 ;
        RECT 54.050 141.435 54.280 141.580 ;
        RECT 54.465 141.505 54.725 141.580 ;
        RECT 55.690 141.435 55.920 141.580 ;
        RECT 57.625 141.435 57.855 141.580 ;
        RECT 58.825 141.435 59.055 141.580 ;
        RECT 59.260 141.550 59.550 142.625 ;
        RECT 60.310 142.625 62.215 142.690 ;
        RECT 64.705 142.625 66.260 142.795 ;
        RECT 67.015 142.795 67.315 143.050 ;
        RECT 67.470 142.935 67.700 143.080 ;
        RECT 69.110 143.005 69.405 143.080 ;
        RECT 69.110 142.935 69.340 143.005 ;
        RECT 71.045 142.935 71.275 143.080 ;
        RECT 72.245 142.935 72.475 143.080 ;
        RECT 67.905 142.795 68.905 142.825 ;
        RECT 71.435 142.795 72.085 142.825 ;
        RECT 72.680 142.795 72.970 144.125 ;
        RECT 73.730 143.050 74.020 145.690 ;
        RECT 74.595 145.625 75.635 145.795 ;
        RECT 78.125 145.625 79.680 145.795 ;
        RECT 80.435 145.690 80.735 146.050 ;
        RECT 80.890 145.935 81.120 146.080 ;
        RECT 81.305 146.005 81.565 146.080 ;
        RECT 82.530 145.935 82.760 146.080 ;
        RECT 84.465 145.935 84.695 146.080 ;
        RECT 85.665 145.935 85.895 146.080 ;
        RECT 81.325 145.795 82.325 145.825 ;
        RECT 84.855 145.795 85.505 145.825 ;
        RECT 86.100 145.795 86.390 146.915 ;
        RECT 87.150 146.050 87.440 146.915 ;
        RECT 88.035 146.705 89.035 146.735 ;
        RECT 90.170 146.705 90.430 146.780 ;
        RECT 91.565 146.705 92.215 146.735 ;
        RECT 88.015 146.535 92.235 146.705 ;
        RECT 88.035 146.505 89.035 146.535 ;
        RECT 90.170 146.460 90.430 146.535 ;
        RECT 91.565 146.505 92.215 146.535 ;
        RECT 87.600 146.250 87.830 146.395 ;
        RECT 88.015 146.250 88.275 146.325 ;
        RECT 89.240 146.250 89.470 146.395 ;
        RECT 91.175 146.250 91.405 146.395 ;
        RECT 92.375 146.250 92.605 146.395 ;
        RECT 87.600 146.080 92.605 146.250 ;
        RECT 74.615 145.595 75.615 145.625 ;
        RECT 78.145 145.595 78.795 145.625 ;
        RECT 75.030 145.235 75.200 145.595 ;
        RECT 74.615 145.205 75.615 145.235 ;
        RECT 76.750 145.205 77.010 145.280 ;
        RECT 78.145 145.205 78.795 145.235 ;
        RECT 74.595 145.035 75.635 145.205 ;
        RECT 76.750 145.035 78.815 145.205 ;
        RECT 74.615 145.005 75.615 145.035 ;
        RECT 76.750 144.960 77.010 145.035 ;
        RECT 78.145 145.005 78.795 145.035 ;
        RECT 74.180 144.750 74.410 144.895 ;
        RECT 75.820 144.825 76.050 144.895 ;
        RECT 75.435 144.750 76.050 144.825 ;
        RECT 77.755 144.750 77.985 144.895 ;
        RECT 78.955 144.750 79.185 144.895 ;
        RECT 74.180 144.580 79.185 144.750 ;
        RECT 74.180 144.435 74.410 144.580 ;
        RECT 75.435 144.505 76.050 144.580 ;
        RECT 75.820 144.435 76.050 144.505 ;
        RECT 77.755 144.435 77.985 144.580 ;
        RECT 78.955 144.435 79.185 144.580 ;
        RECT 79.390 144.550 79.680 145.625 ;
        RECT 74.615 144.295 75.615 144.325 ;
        RECT 78.145 144.295 78.795 144.325 ;
        RECT 79.385 144.295 79.685 144.550 ;
        RECT 74.595 144.125 75.635 144.295 ;
        RECT 78.125 144.190 79.685 144.295 ;
        RECT 78.125 144.125 79.680 144.190 ;
        RECT 74.615 144.095 75.615 144.125 ;
        RECT 78.145 144.095 78.795 144.125 ;
        RECT 75.030 143.735 75.200 144.095 ;
        RECT 74.615 143.705 75.615 143.735 ;
        RECT 76.750 143.705 77.010 143.780 ;
        RECT 78.145 143.705 78.795 143.735 ;
        RECT 74.595 143.535 75.635 143.705 ;
        RECT 76.750 143.535 78.815 143.705 ;
        RECT 74.615 143.505 75.615 143.535 ;
        RECT 76.750 143.460 77.010 143.535 ;
        RECT 78.145 143.505 78.795 143.535 ;
        RECT 74.180 143.250 74.410 143.395 ;
        RECT 75.820 143.325 76.050 143.395 ;
        RECT 75.820 143.250 76.115 143.325 ;
        RECT 77.755 143.250 77.985 143.395 ;
        RECT 78.955 143.250 79.185 143.395 ;
        RECT 74.180 143.080 79.185 143.250 ;
        RECT 67.015 142.690 68.925 142.795 ;
        RECT 54.485 141.295 55.485 141.325 ;
        RECT 58.015 141.295 58.665 141.325 ;
        RECT 59.255 141.295 59.555 141.550 ;
        RECT 54.465 141.125 55.505 141.295 ;
        RECT 57.995 141.190 59.555 141.295 ;
        RECT 57.995 141.125 59.550 141.190 ;
        RECT 54.485 141.095 55.485 141.125 ;
        RECT 58.015 141.095 58.665 141.125 ;
        RECT 54.900 140.735 55.070 141.095 ;
        RECT 54.485 140.705 55.485 140.735 ;
        RECT 56.620 140.705 56.880 140.780 ;
        RECT 58.015 140.705 58.665 140.735 ;
        RECT 54.465 140.535 55.505 140.705 ;
        RECT 56.620 140.535 58.685 140.705 ;
        RECT 54.485 140.505 55.485 140.535 ;
        RECT 56.620 140.460 56.880 140.535 ;
        RECT 58.015 140.505 58.665 140.535 ;
        RECT 54.050 140.250 54.280 140.395 ;
        RECT 54.885 140.250 55.145 140.325 ;
        RECT 55.690 140.250 55.920 140.395 ;
        RECT 57.625 140.250 57.855 140.395 ;
        RECT 58.825 140.250 59.055 140.395 ;
        RECT 54.050 140.080 59.055 140.250 ;
        RECT 41.065 139.595 42.065 139.625 ;
        RECT 44.595 139.595 45.245 139.625 ;
        RECT 41.480 139.235 41.650 139.595 ;
        RECT 41.065 139.205 42.065 139.235 ;
        RECT 43.200 139.205 43.460 139.280 ;
        RECT 44.595 139.205 45.245 139.235 ;
        RECT 41.045 139.035 42.085 139.205 ;
        RECT 43.200 139.035 45.265 139.205 ;
        RECT 41.065 139.005 42.065 139.035 ;
        RECT 43.200 138.960 43.460 139.035 ;
        RECT 44.595 139.005 45.245 139.035 ;
        RECT 40.630 138.750 40.860 138.895 ;
        RECT 42.270 138.825 42.500 138.895 ;
        RECT 42.270 138.750 42.565 138.825 ;
        RECT 44.205 138.750 44.435 138.895 ;
        RECT 45.405 138.750 45.635 138.895 ;
        RECT 40.630 138.580 45.635 138.750 ;
        RECT 40.630 138.435 40.860 138.580 ;
        RECT 42.270 138.505 42.565 138.580 ;
        RECT 42.270 138.435 42.500 138.505 ;
        RECT 44.205 138.435 44.435 138.580 ;
        RECT 45.405 138.435 45.635 138.580 ;
        RECT 45.840 138.550 46.130 139.625 ;
        RECT 41.065 138.295 42.065 138.325 ;
        RECT 44.595 138.295 45.245 138.325 ;
        RECT 45.835 138.295 46.135 138.550 ;
        RECT 37.865 138.125 39.420 138.190 ;
        RECT 33.470 137.050 33.760 138.125 ;
        RECT 34.355 138.095 35.355 138.125 ;
        RECT 37.885 138.095 38.535 138.125 ;
        RECT 34.755 137.735 35.015 137.780 ;
        RECT 34.355 137.705 35.355 137.735 ;
        RECT 37.885 137.705 38.535 137.735 ;
        RECT 34.335 137.535 38.555 137.705 ;
        RECT 34.355 137.505 35.355 137.535 ;
        RECT 37.885 137.505 38.535 137.535 ;
        RECT 34.755 137.460 35.015 137.505 ;
        RECT 33.920 137.250 34.150 137.395 ;
        RECT 35.560 137.250 35.790 137.395 ;
        RECT 36.490 137.250 36.750 137.325 ;
        RECT 37.495 137.250 37.725 137.395 ;
        RECT 38.695 137.250 38.925 137.395 ;
        RECT 33.920 137.080 38.925 137.250 ;
        RECT 26.755 136.690 28.665 136.795 ;
        RECT 26.760 136.625 28.665 136.690 ;
        RECT 26.760 135.295 27.050 136.625 ;
        RECT 27.645 136.595 28.645 136.625 ;
        RECT 28.890 136.365 29.150 136.685 ;
        RECT 31.155 136.625 32.710 136.795 ;
        RECT 33.465 136.795 33.765 137.050 ;
        RECT 33.920 136.935 34.150 137.080 ;
        RECT 35.560 136.935 35.790 137.080 ;
        RECT 36.490 137.005 36.750 137.080 ;
        RECT 37.495 136.935 37.725 137.080 ;
        RECT 38.695 136.935 38.925 137.080 ;
        RECT 34.355 136.795 35.355 136.825 ;
        RECT 37.885 136.795 38.535 136.825 ;
        RECT 39.130 136.795 39.420 138.125 ;
        RECT 40.180 138.125 42.085 138.295 ;
        RECT 44.575 138.190 46.135 138.295 ;
        RECT 46.890 138.295 47.180 139.690 ;
        RECT 47.755 139.625 48.795 139.795 ;
        RECT 51.285 139.625 52.840 139.795 ;
        RECT 53.595 139.690 53.895 140.050 ;
        RECT 54.050 139.935 54.280 140.080 ;
        RECT 54.885 140.005 55.145 140.080 ;
        RECT 55.690 139.935 55.920 140.080 ;
        RECT 57.625 139.935 57.855 140.080 ;
        RECT 58.825 139.935 59.055 140.080 ;
        RECT 54.485 139.795 55.485 139.825 ;
        RECT 58.015 139.795 58.665 139.825 ;
        RECT 59.260 139.795 59.550 141.125 ;
        RECT 60.310 140.050 60.600 142.625 ;
        RECT 61.195 142.595 62.195 142.625 ;
        RECT 64.725 142.595 65.375 142.625 ;
        RECT 61.195 142.205 62.195 142.235 ;
        RECT 63.330 142.205 63.590 142.280 ;
        RECT 64.725 142.205 65.375 142.235 ;
        RECT 61.175 142.035 65.395 142.205 ;
        RECT 61.195 142.005 62.195 142.035 ;
        RECT 63.330 141.960 63.590 142.035 ;
        RECT 64.725 142.005 65.375 142.035 ;
        RECT 60.760 141.750 60.990 141.895 ;
        RECT 61.175 141.750 61.435 141.825 ;
        RECT 62.400 141.750 62.630 141.895 ;
        RECT 64.335 141.750 64.565 141.895 ;
        RECT 65.535 141.750 65.765 141.895 ;
        RECT 60.760 141.580 65.765 141.750 ;
        RECT 60.760 141.435 60.990 141.580 ;
        RECT 61.175 141.505 61.435 141.580 ;
        RECT 62.400 141.435 62.630 141.580 ;
        RECT 64.335 141.435 64.565 141.580 ;
        RECT 65.535 141.435 65.765 141.580 ;
        RECT 65.970 141.550 66.260 142.625 ;
        RECT 67.020 142.625 68.925 142.690 ;
        RECT 71.415 142.625 72.970 142.795 ;
        RECT 73.725 142.795 74.025 143.050 ;
        RECT 74.180 142.935 74.410 143.080 ;
        RECT 75.820 143.005 76.115 143.080 ;
        RECT 75.820 142.935 76.050 143.005 ;
        RECT 77.755 142.935 77.985 143.080 ;
        RECT 78.955 142.935 79.185 143.080 ;
        RECT 74.615 142.795 75.615 142.825 ;
        RECT 78.145 142.795 78.795 142.825 ;
        RECT 79.390 142.795 79.680 144.125 ;
        RECT 80.440 143.050 80.730 145.690 ;
        RECT 81.305 145.625 82.345 145.795 ;
        RECT 84.835 145.625 86.390 145.795 ;
        RECT 87.145 145.690 87.445 146.050 ;
        RECT 87.600 145.935 87.830 146.080 ;
        RECT 88.015 146.005 88.275 146.080 ;
        RECT 89.240 145.935 89.470 146.080 ;
        RECT 91.175 145.935 91.405 146.080 ;
        RECT 92.375 145.935 92.605 146.080 ;
        RECT 88.035 145.795 89.035 145.825 ;
        RECT 91.565 145.795 92.215 145.825 ;
        RECT 92.810 145.795 93.100 146.915 ;
        RECT 81.325 145.595 82.325 145.625 ;
        RECT 84.855 145.595 85.505 145.625 ;
        RECT 81.740 145.235 81.910 145.595 ;
        RECT 81.325 145.205 82.325 145.235 ;
        RECT 83.460 145.205 83.720 145.280 ;
        RECT 84.855 145.205 85.505 145.235 ;
        RECT 81.305 145.035 82.345 145.205 ;
        RECT 83.460 145.035 85.525 145.205 ;
        RECT 81.325 145.005 82.325 145.035 ;
        RECT 83.460 144.960 83.720 145.035 ;
        RECT 84.855 145.005 85.505 145.035 ;
        RECT 80.890 144.750 81.120 144.895 ;
        RECT 82.530 144.825 82.760 144.895 ;
        RECT 82.145 144.750 82.760 144.825 ;
        RECT 84.465 144.750 84.695 144.895 ;
        RECT 85.665 144.750 85.895 144.895 ;
        RECT 80.890 144.580 85.895 144.750 ;
        RECT 80.890 144.435 81.120 144.580 ;
        RECT 82.145 144.505 82.760 144.580 ;
        RECT 82.530 144.435 82.760 144.505 ;
        RECT 84.465 144.435 84.695 144.580 ;
        RECT 85.665 144.435 85.895 144.580 ;
        RECT 86.100 144.550 86.390 145.625 ;
        RECT 81.325 144.295 82.325 144.325 ;
        RECT 84.855 144.295 85.505 144.325 ;
        RECT 86.095 144.295 86.395 144.550 ;
        RECT 81.305 144.125 82.345 144.295 ;
        RECT 84.835 144.190 86.395 144.295 ;
        RECT 84.835 144.125 86.390 144.190 ;
        RECT 81.325 144.095 82.325 144.125 ;
        RECT 84.855 144.095 85.505 144.125 ;
        RECT 81.740 143.735 81.910 144.095 ;
        RECT 81.325 143.705 82.325 143.735 ;
        RECT 83.460 143.705 83.720 143.780 ;
        RECT 84.855 143.705 85.505 143.735 ;
        RECT 81.305 143.535 82.345 143.705 ;
        RECT 83.460 143.535 85.525 143.705 ;
        RECT 81.325 143.505 82.325 143.535 ;
        RECT 83.460 143.460 83.720 143.535 ;
        RECT 84.855 143.505 85.505 143.535 ;
        RECT 80.890 143.250 81.120 143.395 ;
        RECT 82.530 143.325 82.760 143.395 ;
        RECT 82.530 143.250 82.825 143.325 ;
        RECT 84.465 143.250 84.695 143.395 ;
        RECT 85.665 143.250 85.895 143.395 ;
        RECT 80.890 143.080 85.895 143.250 ;
        RECT 73.725 142.690 75.635 142.795 ;
        RECT 61.195 141.295 62.195 141.325 ;
        RECT 64.725 141.295 65.375 141.325 ;
        RECT 65.965 141.295 66.265 141.550 ;
        RECT 61.175 141.125 62.215 141.295 ;
        RECT 64.705 141.190 66.265 141.295 ;
        RECT 64.705 141.125 66.260 141.190 ;
        RECT 61.195 141.095 62.195 141.125 ;
        RECT 64.725 141.095 65.375 141.125 ;
        RECT 61.610 140.735 61.780 141.095 ;
        RECT 61.195 140.705 62.195 140.735 ;
        RECT 63.330 140.705 63.590 140.780 ;
        RECT 64.725 140.705 65.375 140.735 ;
        RECT 61.175 140.535 62.215 140.705 ;
        RECT 63.330 140.535 65.395 140.705 ;
        RECT 61.195 140.505 62.195 140.535 ;
        RECT 63.330 140.460 63.590 140.535 ;
        RECT 64.725 140.505 65.375 140.535 ;
        RECT 60.760 140.250 60.990 140.395 ;
        RECT 61.595 140.250 61.855 140.325 ;
        RECT 62.400 140.250 62.630 140.395 ;
        RECT 64.335 140.250 64.565 140.395 ;
        RECT 65.535 140.250 65.765 140.395 ;
        RECT 60.760 140.080 65.765 140.250 ;
        RECT 47.775 139.595 48.775 139.625 ;
        RECT 51.305 139.595 51.955 139.625 ;
        RECT 48.190 139.235 48.360 139.595 ;
        RECT 47.775 139.205 48.775 139.235 ;
        RECT 49.910 139.205 50.170 139.280 ;
        RECT 51.305 139.205 51.955 139.235 ;
        RECT 47.755 139.035 48.795 139.205 ;
        RECT 49.910 139.035 51.975 139.205 ;
        RECT 47.775 139.005 48.775 139.035 ;
        RECT 49.910 138.960 50.170 139.035 ;
        RECT 51.305 139.005 51.955 139.035 ;
        RECT 47.340 138.750 47.570 138.895 ;
        RECT 48.980 138.825 49.210 138.895 ;
        RECT 48.980 138.750 49.275 138.825 ;
        RECT 50.915 138.750 51.145 138.895 ;
        RECT 52.115 138.750 52.345 138.895 ;
        RECT 47.340 138.580 52.345 138.750 ;
        RECT 47.340 138.435 47.570 138.580 ;
        RECT 48.980 138.505 49.275 138.580 ;
        RECT 48.980 138.435 49.210 138.505 ;
        RECT 50.915 138.435 51.145 138.580 ;
        RECT 52.115 138.435 52.345 138.580 ;
        RECT 52.550 138.550 52.840 139.625 ;
        RECT 47.775 138.295 48.775 138.325 ;
        RECT 51.305 138.295 51.955 138.325 ;
        RECT 52.545 138.295 52.845 138.550 ;
        RECT 44.575 138.125 46.130 138.190 ;
        RECT 40.180 137.050 40.470 138.125 ;
        RECT 41.065 138.095 42.065 138.125 ;
        RECT 44.595 138.095 45.245 138.125 ;
        RECT 45.005 137.735 45.265 137.780 ;
        RECT 41.065 137.705 42.065 137.735 ;
        RECT 44.595 137.705 45.265 137.735 ;
        RECT 41.045 137.535 45.265 137.705 ;
        RECT 41.065 137.505 42.065 137.535 ;
        RECT 44.595 137.505 45.265 137.535 ;
        RECT 45.005 137.460 45.265 137.505 ;
        RECT 40.630 137.250 40.860 137.395 ;
        RECT 42.270 137.250 42.500 137.395 ;
        RECT 43.200 137.250 43.460 137.325 ;
        RECT 44.205 137.250 44.435 137.395 ;
        RECT 45.405 137.250 45.635 137.395 ;
        RECT 40.630 137.080 45.635 137.250 ;
        RECT 33.465 136.690 35.375 136.795 ;
        RECT 31.175 136.595 31.825 136.625 ;
        RECT 27.645 136.205 28.645 136.235 ;
        RECT 28.935 136.205 29.105 136.365 ;
        RECT 29.780 136.205 30.040 136.280 ;
        RECT 31.175 136.205 31.825 136.235 ;
        RECT 27.625 136.035 31.845 136.205 ;
        RECT 27.645 136.005 28.645 136.035 ;
        RECT 29.780 135.960 30.040 136.035 ;
        RECT 31.175 136.005 31.825 136.035 ;
        RECT 27.210 135.750 27.440 135.895 ;
        RECT 28.850 135.750 29.080 135.895 ;
        RECT 29.750 135.750 30.070 135.795 ;
        RECT 30.785 135.750 31.015 135.895 ;
        RECT 31.985 135.750 32.215 135.895 ;
        RECT 27.210 135.580 32.215 135.750 ;
        RECT 27.210 135.435 27.440 135.580 ;
        RECT 28.850 135.435 29.080 135.580 ;
        RECT 29.750 135.535 30.070 135.580 ;
        RECT 30.785 135.435 31.015 135.580 ;
        RECT 31.985 135.435 32.215 135.580 ;
        RECT 32.420 135.550 32.710 136.625 ;
        RECT 33.470 136.625 35.375 136.690 ;
        RECT 37.865 136.625 39.420 136.795 ;
        RECT 40.175 136.795 40.475 137.050 ;
        RECT 40.630 136.935 40.860 137.080 ;
        RECT 42.270 136.935 42.500 137.080 ;
        RECT 43.200 137.005 43.460 137.080 ;
        RECT 44.205 136.935 44.435 137.080 ;
        RECT 45.405 136.935 45.635 137.080 ;
        RECT 41.065 136.795 42.065 136.825 ;
        RECT 44.595 136.795 45.245 136.825 ;
        RECT 45.840 136.795 46.130 138.125 ;
        RECT 46.890 138.125 48.795 138.295 ;
        RECT 51.285 138.190 52.845 138.295 ;
        RECT 53.600 138.295 53.890 139.690 ;
        RECT 54.465 139.625 55.505 139.795 ;
        RECT 57.995 139.625 59.550 139.795 ;
        RECT 60.305 139.690 60.605 140.050 ;
        RECT 60.760 139.935 60.990 140.080 ;
        RECT 61.595 140.005 61.855 140.080 ;
        RECT 62.400 139.935 62.630 140.080 ;
        RECT 64.335 139.935 64.565 140.080 ;
        RECT 65.535 139.935 65.765 140.080 ;
        RECT 61.195 139.795 62.195 139.825 ;
        RECT 64.725 139.795 65.375 139.825 ;
        RECT 65.970 139.795 66.260 141.125 ;
        RECT 67.020 140.050 67.310 142.625 ;
        RECT 67.905 142.595 68.905 142.625 ;
        RECT 71.435 142.595 72.085 142.625 ;
        RECT 67.905 142.205 68.905 142.235 ;
        RECT 70.040 142.205 70.300 142.280 ;
        RECT 71.435 142.205 72.085 142.235 ;
        RECT 67.885 142.035 72.105 142.205 ;
        RECT 67.905 142.005 68.905 142.035 ;
        RECT 70.040 141.960 70.300 142.035 ;
        RECT 71.435 142.005 72.085 142.035 ;
        RECT 67.470 141.750 67.700 141.895 ;
        RECT 67.885 141.750 68.145 141.825 ;
        RECT 69.110 141.750 69.340 141.895 ;
        RECT 71.045 141.750 71.275 141.895 ;
        RECT 72.245 141.750 72.475 141.895 ;
        RECT 67.470 141.580 72.475 141.750 ;
        RECT 67.470 141.435 67.700 141.580 ;
        RECT 67.885 141.505 68.145 141.580 ;
        RECT 69.110 141.435 69.340 141.580 ;
        RECT 71.045 141.435 71.275 141.580 ;
        RECT 72.245 141.435 72.475 141.580 ;
        RECT 72.680 141.550 72.970 142.625 ;
        RECT 73.730 142.625 75.635 142.690 ;
        RECT 78.125 142.625 79.680 142.795 ;
        RECT 80.435 142.795 80.735 143.050 ;
        RECT 80.890 142.935 81.120 143.080 ;
        RECT 82.530 143.005 82.825 143.080 ;
        RECT 82.530 142.935 82.760 143.005 ;
        RECT 84.465 142.935 84.695 143.080 ;
        RECT 85.665 142.935 85.895 143.080 ;
        RECT 81.325 142.795 82.325 142.825 ;
        RECT 84.855 142.795 85.505 142.825 ;
        RECT 86.100 142.795 86.390 144.125 ;
        RECT 87.150 143.050 87.440 145.690 ;
        RECT 88.015 145.625 89.055 145.795 ;
        RECT 91.545 145.625 93.100 145.795 ;
        RECT 88.035 145.595 89.035 145.625 ;
        RECT 91.565 145.595 92.215 145.625 ;
        RECT 88.450 145.235 88.620 145.595 ;
        RECT 88.035 145.205 89.035 145.235 ;
        RECT 90.170 145.205 90.430 145.280 ;
        RECT 91.565 145.205 92.215 145.235 ;
        RECT 88.015 145.035 89.055 145.205 ;
        RECT 90.170 145.035 92.235 145.205 ;
        RECT 88.035 145.005 89.035 145.035 ;
        RECT 90.170 144.960 90.430 145.035 ;
        RECT 91.565 145.005 92.215 145.035 ;
        RECT 87.600 144.750 87.830 144.895 ;
        RECT 89.240 144.825 89.470 144.895 ;
        RECT 88.855 144.750 89.470 144.825 ;
        RECT 91.175 144.750 91.405 144.895 ;
        RECT 92.375 144.750 92.605 144.895 ;
        RECT 87.600 144.580 92.605 144.750 ;
        RECT 87.600 144.435 87.830 144.580 ;
        RECT 88.855 144.505 89.470 144.580 ;
        RECT 89.240 144.435 89.470 144.505 ;
        RECT 91.175 144.435 91.405 144.580 ;
        RECT 92.375 144.435 92.605 144.580 ;
        RECT 92.810 144.550 93.100 145.625 ;
        RECT 88.035 144.295 89.035 144.325 ;
        RECT 91.565 144.295 92.215 144.325 ;
        RECT 92.805 144.295 93.105 144.550 ;
        RECT 88.015 144.125 89.055 144.295 ;
        RECT 91.545 144.190 93.105 144.295 ;
        RECT 91.545 144.125 93.100 144.190 ;
        RECT 88.035 144.095 89.035 144.125 ;
        RECT 91.565 144.095 92.215 144.125 ;
        RECT 88.450 143.735 88.620 144.095 ;
        RECT 88.035 143.705 89.035 143.735 ;
        RECT 90.170 143.705 90.430 143.780 ;
        RECT 91.565 143.705 92.215 143.735 ;
        RECT 88.015 143.535 89.055 143.705 ;
        RECT 90.170 143.535 92.235 143.705 ;
        RECT 88.035 143.505 89.035 143.535 ;
        RECT 90.170 143.460 90.430 143.535 ;
        RECT 91.565 143.505 92.215 143.535 ;
        RECT 87.600 143.250 87.830 143.395 ;
        RECT 89.240 143.325 89.470 143.395 ;
        RECT 89.240 143.250 89.535 143.325 ;
        RECT 91.175 143.250 91.405 143.395 ;
        RECT 92.375 143.250 92.605 143.395 ;
        RECT 87.600 143.080 92.605 143.250 ;
        RECT 80.435 142.690 82.345 142.795 ;
        RECT 67.905 141.295 68.905 141.325 ;
        RECT 71.435 141.295 72.085 141.325 ;
        RECT 72.675 141.295 72.975 141.550 ;
        RECT 67.885 141.125 68.925 141.295 ;
        RECT 71.415 141.190 72.975 141.295 ;
        RECT 71.415 141.125 72.970 141.190 ;
        RECT 67.905 141.095 68.905 141.125 ;
        RECT 71.435 141.095 72.085 141.125 ;
        RECT 68.320 140.735 68.490 141.095 ;
        RECT 67.905 140.705 68.905 140.735 ;
        RECT 70.040 140.705 70.300 140.780 ;
        RECT 71.435 140.705 72.085 140.735 ;
        RECT 67.885 140.535 68.925 140.705 ;
        RECT 70.040 140.535 72.105 140.705 ;
        RECT 67.905 140.505 68.905 140.535 ;
        RECT 70.040 140.460 70.300 140.535 ;
        RECT 71.435 140.505 72.085 140.535 ;
        RECT 67.470 140.250 67.700 140.395 ;
        RECT 68.305 140.250 68.565 140.325 ;
        RECT 69.110 140.250 69.340 140.395 ;
        RECT 71.045 140.250 71.275 140.395 ;
        RECT 72.245 140.250 72.475 140.395 ;
        RECT 67.470 140.080 72.475 140.250 ;
        RECT 54.485 139.595 55.485 139.625 ;
        RECT 58.015 139.595 58.665 139.625 ;
        RECT 54.900 139.235 55.070 139.595 ;
        RECT 54.485 139.205 55.485 139.235 ;
        RECT 56.620 139.205 56.880 139.280 ;
        RECT 58.015 139.205 58.665 139.235 ;
        RECT 54.465 139.035 55.505 139.205 ;
        RECT 56.620 139.035 58.685 139.205 ;
        RECT 54.485 139.005 55.485 139.035 ;
        RECT 56.620 138.960 56.880 139.035 ;
        RECT 58.015 139.005 58.665 139.035 ;
        RECT 54.050 138.750 54.280 138.895 ;
        RECT 55.690 138.825 55.920 138.895 ;
        RECT 55.690 138.750 55.985 138.825 ;
        RECT 57.625 138.750 57.855 138.895 ;
        RECT 58.825 138.750 59.055 138.895 ;
        RECT 54.050 138.580 59.055 138.750 ;
        RECT 54.050 138.435 54.280 138.580 ;
        RECT 55.690 138.505 55.985 138.580 ;
        RECT 55.690 138.435 55.920 138.505 ;
        RECT 57.625 138.435 57.855 138.580 ;
        RECT 58.825 138.435 59.055 138.580 ;
        RECT 59.260 138.550 59.550 139.625 ;
        RECT 54.485 138.295 55.485 138.325 ;
        RECT 58.015 138.295 58.665 138.325 ;
        RECT 59.255 138.295 59.555 138.550 ;
        RECT 51.285 138.125 52.840 138.190 ;
        RECT 46.890 137.050 47.180 138.125 ;
        RECT 47.775 138.095 48.775 138.125 ;
        RECT 51.305 138.095 51.955 138.125 ;
        RECT 48.175 137.735 48.435 137.780 ;
        RECT 47.775 137.705 48.775 137.735 ;
        RECT 51.305 137.705 51.955 137.735 ;
        RECT 47.755 137.535 51.975 137.705 ;
        RECT 47.775 137.505 48.775 137.535 ;
        RECT 51.305 137.505 51.955 137.535 ;
        RECT 48.175 137.460 48.435 137.505 ;
        RECT 47.340 137.250 47.570 137.395 ;
        RECT 48.980 137.250 49.210 137.395 ;
        RECT 49.910 137.250 50.170 137.325 ;
        RECT 50.915 137.250 51.145 137.395 ;
        RECT 52.115 137.250 52.345 137.395 ;
        RECT 47.340 137.080 52.345 137.250 ;
        RECT 40.175 136.690 42.085 136.795 ;
        RECT 27.645 135.295 28.645 135.325 ;
        RECT 31.175 135.295 31.825 135.325 ;
        RECT 32.415 135.295 32.715 135.550 ;
        RECT 26.760 135.125 28.665 135.295 ;
        RECT 31.155 135.190 32.715 135.295 ;
        RECT 33.470 135.295 33.760 136.625 ;
        RECT 34.355 136.595 35.355 136.625 ;
        RECT 37.885 136.595 38.535 136.625 ;
        RECT 35.175 136.235 35.435 136.280 ;
        RECT 34.355 136.205 35.435 136.235 ;
        RECT 36.490 136.205 36.750 136.280 ;
        RECT 37.885 136.205 38.535 136.235 ;
        RECT 34.335 136.035 38.555 136.205 ;
        RECT 34.355 136.005 35.435 136.035 ;
        RECT 35.175 135.960 35.435 136.005 ;
        RECT 36.490 135.960 36.750 136.035 ;
        RECT 37.885 136.005 38.535 136.035 ;
        RECT 33.920 135.750 34.150 135.895 ;
        RECT 35.560 135.750 35.790 135.895 ;
        RECT 36.460 135.750 36.780 135.795 ;
        RECT 37.495 135.750 37.725 135.895 ;
        RECT 38.695 135.750 38.925 135.895 ;
        RECT 33.920 135.580 38.925 135.750 ;
        RECT 33.920 135.435 34.150 135.580 ;
        RECT 35.560 135.435 35.790 135.580 ;
        RECT 36.460 135.535 36.780 135.580 ;
        RECT 37.495 135.435 37.725 135.580 ;
        RECT 38.695 135.435 38.925 135.580 ;
        RECT 39.130 135.550 39.420 136.625 ;
        RECT 40.180 136.625 42.085 136.690 ;
        RECT 34.355 135.295 35.355 135.325 ;
        RECT 37.885 135.295 38.535 135.325 ;
        RECT 39.125 135.295 39.425 135.550 ;
        RECT 31.155 135.125 32.710 135.190 ;
        RECT 26.760 134.050 27.050 135.125 ;
        RECT 27.645 135.095 28.645 135.125 ;
        RECT 31.175 135.095 31.825 135.125 ;
        RECT 27.645 134.705 28.645 134.735 ;
        RECT 31.175 134.705 31.825 134.735 ;
        RECT 27.625 134.535 31.845 134.705 ;
        RECT 27.645 134.505 28.645 134.535 ;
        RECT 31.175 134.505 31.825 134.535 ;
        RECT 27.210 134.250 27.440 134.395 ;
        RECT 28.850 134.250 29.080 134.395 ;
        RECT 30.785 134.250 31.015 134.395 ;
        RECT 31.985 134.250 32.215 134.395 ;
        RECT 32.420 134.250 32.710 135.125 ;
        RECT 27.210 134.080 32.710 134.250 ;
        RECT 26.755 133.795 27.055 134.050 ;
        RECT 27.210 133.935 27.440 134.080 ;
        RECT 28.850 133.935 29.080 134.080 ;
        RECT 30.785 133.935 31.015 134.080 ;
        RECT 31.985 133.935 32.215 134.080 ;
        RECT 27.645 133.795 28.645 133.825 ;
        RECT 31.175 133.795 31.825 133.825 ;
        RECT 32.420 133.795 32.710 134.080 ;
        RECT 33.470 135.125 35.375 135.295 ;
        RECT 37.865 135.190 39.425 135.295 ;
        RECT 40.180 135.295 40.470 136.625 ;
        RECT 41.065 136.595 42.065 136.625 ;
        RECT 42.310 136.365 42.570 136.685 ;
        RECT 44.575 136.625 46.130 136.795 ;
        RECT 46.885 136.795 47.185 137.050 ;
        RECT 47.340 136.935 47.570 137.080 ;
        RECT 48.980 136.935 49.210 137.080 ;
        RECT 49.910 137.005 50.170 137.080 ;
        RECT 50.915 136.935 51.145 137.080 ;
        RECT 52.115 136.935 52.345 137.080 ;
        RECT 47.775 136.795 48.775 136.825 ;
        RECT 51.305 136.795 51.955 136.825 ;
        RECT 52.550 136.795 52.840 138.125 ;
        RECT 53.600 138.125 55.505 138.295 ;
        RECT 57.995 138.190 59.555 138.295 ;
        RECT 60.310 138.295 60.600 139.690 ;
        RECT 61.175 139.625 62.215 139.795 ;
        RECT 64.705 139.625 66.260 139.795 ;
        RECT 67.015 139.690 67.315 140.050 ;
        RECT 67.470 139.935 67.700 140.080 ;
        RECT 68.305 140.005 68.565 140.080 ;
        RECT 69.110 139.935 69.340 140.080 ;
        RECT 71.045 139.935 71.275 140.080 ;
        RECT 72.245 139.935 72.475 140.080 ;
        RECT 67.905 139.795 68.905 139.825 ;
        RECT 71.435 139.795 72.085 139.825 ;
        RECT 72.680 139.795 72.970 141.125 ;
        RECT 73.730 140.050 74.020 142.625 ;
        RECT 74.615 142.595 75.615 142.625 ;
        RECT 78.145 142.595 78.795 142.625 ;
        RECT 74.615 142.205 75.615 142.235 ;
        RECT 76.750 142.205 77.010 142.280 ;
        RECT 78.145 142.205 78.795 142.235 ;
        RECT 74.595 142.035 78.815 142.205 ;
        RECT 74.615 142.005 75.615 142.035 ;
        RECT 76.750 141.960 77.010 142.035 ;
        RECT 78.145 142.005 78.795 142.035 ;
        RECT 74.180 141.750 74.410 141.895 ;
        RECT 74.595 141.750 74.855 141.825 ;
        RECT 75.820 141.750 76.050 141.895 ;
        RECT 77.755 141.750 77.985 141.895 ;
        RECT 78.955 141.750 79.185 141.895 ;
        RECT 74.180 141.580 79.185 141.750 ;
        RECT 74.180 141.435 74.410 141.580 ;
        RECT 74.595 141.505 74.855 141.580 ;
        RECT 75.820 141.435 76.050 141.580 ;
        RECT 77.755 141.435 77.985 141.580 ;
        RECT 78.955 141.435 79.185 141.580 ;
        RECT 79.390 141.550 79.680 142.625 ;
        RECT 80.440 142.625 82.345 142.690 ;
        RECT 84.835 142.625 86.390 142.795 ;
        RECT 87.145 142.795 87.445 143.050 ;
        RECT 87.600 142.935 87.830 143.080 ;
        RECT 89.240 143.005 89.535 143.080 ;
        RECT 89.240 142.935 89.470 143.005 ;
        RECT 91.175 142.935 91.405 143.080 ;
        RECT 92.375 142.935 92.605 143.080 ;
        RECT 88.035 142.795 89.035 142.825 ;
        RECT 91.565 142.795 92.215 142.825 ;
        RECT 92.810 142.795 93.100 144.125 ;
        RECT 87.145 142.690 89.055 142.795 ;
        RECT 74.615 141.295 75.615 141.325 ;
        RECT 78.145 141.295 78.795 141.325 ;
        RECT 79.385 141.295 79.685 141.550 ;
        RECT 74.595 141.125 75.635 141.295 ;
        RECT 78.125 141.190 79.685 141.295 ;
        RECT 78.125 141.125 79.680 141.190 ;
        RECT 74.615 141.095 75.615 141.125 ;
        RECT 78.145 141.095 78.795 141.125 ;
        RECT 75.030 140.735 75.200 141.095 ;
        RECT 74.615 140.705 75.615 140.735 ;
        RECT 76.750 140.705 77.010 140.780 ;
        RECT 78.145 140.705 78.795 140.735 ;
        RECT 74.595 140.535 75.635 140.705 ;
        RECT 76.750 140.535 78.815 140.705 ;
        RECT 74.615 140.505 75.615 140.535 ;
        RECT 76.750 140.460 77.010 140.535 ;
        RECT 78.145 140.505 78.795 140.535 ;
        RECT 74.180 140.250 74.410 140.395 ;
        RECT 75.015 140.250 75.275 140.325 ;
        RECT 75.820 140.250 76.050 140.395 ;
        RECT 77.755 140.250 77.985 140.395 ;
        RECT 78.955 140.250 79.185 140.395 ;
        RECT 74.180 140.080 79.185 140.250 ;
        RECT 61.195 139.595 62.195 139.625 ;
        RECT 64.725 139.595 65.375 139.625 ;
        RECT 61.610 139.235 61.780 139.595 ;
        RECT 61.195 139.205 62.195 139.235 ;
        RECT 63.330 139.205 63.590 139.280 ;
        RECT 64.725 139.205 65.375 139.235 ;
        RECT 61.175 139.035 62.215 139.205 ;
        RECT 63.330 139.035 65.395 139.205 ;
        RECT 61.195 139.005 62.195 139.035 ;
        RECT 63.330 138.960 63.590 139.035 ;
        RECT 64.725 139.005 65.375 139.035 ;
        RECT 60.760 138.750 60.990 138.895 ;
        RECT 62.400 138.825 62.630 138.895 ;
        RECT 62.400 138.750 62.695 138.825 ;
        RECT 64.335 138.750 64.565 138.895 ;
        RECT 65.535 138.750 65.765 138.895 ;
        RECT 60.760 138.580 65.765 138.750 ;
        RECT 60.760 138.435 60.990 138.580 ;
        RECT 62.400 138.505 62.695 138.580 ;
        RECT 62.400 138.435 62.630 138.505 ;
        RECT 64.335 138.435 64.565 138.580 ;
        RECT 65.535 138.435 65.765 138.580 ;
        RECT 65.970 138.550 66.260 139.625 ;
        RECT 61.195 138.295 62.195 138.325 ;
        RECT 64.725 138.295 65.375 138.325 ;
        RECT 65.965 138.295 66.265 138.550 ;
        RECT 57.995 138.125 59.550 138.190 ;
        RECT 53.600 137.050 53.890 138.125 ;
        RECT 54.485 138.095 55.485 138.125 ;
        RECT 58.015 138.095 58.665 138.125 ;
        RECT 58.425 137.735 58.685 137.780 ;
        RECT 54.485 137.705 55.485 137.735 ;
        RECT 58.015 137.705 58.685 137.735 ;
        RECT 54.465 137.535 58.685 137.705 ;
        RECT 54.485 137.505 55.485 137.535 ;
        RECT 58.015 137.505 58.685 137.535 ;
        RECT 58.425 137.460 58.685 137.505 ;
        RECT 54.050 137.250 54.280 137.395 ;
        RECT 55.690 137.250 55.920 137.395 ;
        RECT 56.620 137.250 56.880 137.325 ;
        RECT 57.625 137.250 57.855 137.395 ;
        RECT 58.825 137.250 59.055 137.395 ;
        RECT 54.050 137.080 59.055 137.250 ;
        RECT 46.885 136.690 48.795 136.795 ;
        RECT 44.595 136.595 45.245 136.625 ;
        RECT 41.065 136.205 42.065 136.235 ;
        RECT 42.355 136.205 42.525 136.365 ;
        RECT 43.200 136.205 43.460 136.280 ;
        RECT 44.595 136.205 45.245 136.235 ;
        RECT 41.045 136.035 45.265 136.205 ;
        RECT 41.065 136.005 42.065 136.035 ;
        RECT 43.200 135.960 43.460 136.035 ;
        RECT 44.595 136.005 45.245 136.035 ;
        RECT 40.630 135.750 40.860 135.895 ;
        RECT 42.270 135.750 42.500 135.895 ;
        RECT 43.170 135.750 43.490 135.795 ;
        RECT 44.205 135.750 44.435 135.895 ;
        RECT 45.405 135.750 45.635 135.895 ;
        RECT 40.630 135.580 45.635 135.750 ;
        RECT 40.630 135.435 40.860 135.580 ;
        RECT 42.270 135.435 42.500 135.580 ;
        RECT 43.170 135.535 43.490 135.580 ;
        RECT 44.205 135.435 44.435 135.580 ;
        RECT 45.405 135.435 45.635 135.580 ;
        RECT 45.840 135.550 46.130 136.625 ;
        RECT 46.890 136.625 48.795 136.690 ;
        RECT 51.285 136.625 52.840 136.795 ;
        RECT 53.595 136.795 53.895 137.050 ;
        RECT 54.050 136.935 54.280 137.080 ;
        RECT 55.690 136.935 55.920 137.080 ;
        RECT 56.620 137.005 56.880 137.080 ;
        RECT 57.625 136.935 57.855 137.080 ;
        RECT 58.825 136.935 59.055 137.080 ;
        RECT 54.485 136.795 55.485 136.825 ;
        RECT 58.015 136.795 58.665 136.825 ;
        RECT 59.260 136.795 59.550 138.125 ;
        RECT 60.310 138.125 62.215 138.295 ;
        RECT 64.705 138.190 66.265 138.295 ;
        RECT 67.020 138.295 67.310 139.690 ;
        RECT 67.885 139.625 68.925 139.795 ;
        RECT 71.415 139.625 72.970 139.795 ;
        RECT 73.725 139.690 74.025 140.050 ;
        RECT 74.180 139.935 74.410 140.080 ;
        RECT 75.015 140.005 75.275 140.080 ;
        RECT 75.820 139.935 76.050 140.080 ;
        RECT 77.755 139.935 77.985 140.080 ;
        RECT 78.955 139.935 79.185 140.080 ;
        RECT 74.615 139.795 75.615 139.825 ;
        RECT 78.145 139.795 78.795 139.825 ;
        RECT 79.390 139.795 79.680 141.125 ;
        RECT 80.440 140.050 80.730 142.625 ;
        RECT 81.325 142.595 82.325 142.625 ;
        RECT 84.855 142.595 85.505 142.625 ;
        RECT 81.325 142.205 82.325 142.235 ;
        RECT 83.460 142.205 83.720 142.280 ;
        RECT 84.855 142.205 85.505 142.235 ;
        RECT 81.305 142.035 85.525 142.205 ;
        RECT 81.325 142.005 82.325 142.035 ;
        RECT 83.460 141.960 83.720 142.035 ;
        RECT 84.855 142.005 85.505 142.035 ;
        RECT 80.890 141.750 81.120 141.895 ;
        RECT 81.305 141.750 81.565 141.825 ;
        RECT 82.530 141.750 82.760 141.895 ;
        RECT 84.465 141.750 84.695 141.895 ;
        RECT 85.665 141.750 85.895 141.895 ;
        RECT 80.890 141.580 85.895 141.750 ;
        RECT 80.890 141.435 81.120 141.580 ;
        RECT 81.305 141.505 81.565 141.580 ;
        RECT 82.530 141.435 82.760 141.580 ;
        RECT 84.465 141.435 84.695 141.580 ;
        RECT 85.665 141.435 85.895 141.580 ;
        RECT 86.100 141.550 86.390 142.625 ;
        RECT 87.150 142.625 89.055 142.690 ;
        RECT 91.545 142.625 93.100 142.795 ;
        RECT 81.325 141.295 82.325 141.325 ;
        RECT 84.855 141.295 85.505 141.325 ;
        RECT 86.095 141.295 86.395 141.550 ;
        RECT 81.305 141.125 82.345 141.295 ;
        RECT 84.835 141.190 86.395 141.295 ;
        RECT 84.835 141.125 86.390 141.190 ;
        RECT 81.325 141.095 82.325 141.125 ;
        RECT 84.855 141.095 85.505 141.125 ;
        RECT 81.740 140.735 81.910 141.095 ;
        RECT 81.325 140.705 82.325 140.735 ;
        RECT 83.460 140.705 83.720 140.780 ;
        RECT 84.855 140.705 85.505 140.735 ;
        RECT 81.305 140.535 82.345 140.705 ;
        RECT 83.460 140.535 85.525 140.705 ;
        RECT 81.325 140.505 82.325 140.535 ;
        RECT 83.460 140.460 83.720 140.535 ;
        RECT 84.855 140.505 85.505 140.535 ;
        RECT 80.890 140.250 81.120 140.395 ;
        RECT 81.725 140.250 81.985 140.325 ;
        RECT 82.530 140.250 82.760 140.395 ;
        RECT 84.465 140.250 84.695 140.395 ;
        RECT 85.665 140.250 85.895 140.395 ;
        RECT 80.890 140.080 85.895 140.250 ;
        RECT 67.905 139.595 68.905 139.625 ;
        RECT 71.435 139.595 72.085 139.625 ;
        RECT 68.320 139.235 68.490 139.595 ;
        RECT 67.905 139.205 68.905 139.235 ;
        RECT 70.040 139.205 70.300 139.280 ;
        RECT 71.435 139.205 72.085 139.235 ;
        RECT 67.885 139.035 68.925 139.205 ;
        RECT 70.040 139.035 72.105 139.205 ;
        RECT 67.905 139.005 68.905 139.035 ;
        RECT 70.040 138.960 70.300 139.035 ;
        RECT 71.435 139.005 72.085 139.035 ;
        RECT 67.470 138.750 67.700 138.895 ;
        RECT 69.110 138.825 69.340 138.895 ;
        RECT 69.110 138.750 69.405 138.825 ;
        RECT 71.045 138.750 71.275 138.895 ;
        RECT 72.245 138.750 72.475 138.895 ;
        RECT 67.470 138.580 72.475 138.750 ;
        RECT 67.470 138.435 67.700 138.580 ;
        RECT 69.110 138.505 69.405 138.580 ;
        RECT 69.110 138.435 69.340 138.505 ;
        RECT 71.045 138.435 71.275 138.580 ;
        RECT 72.245 138.435 72.475 138.580 ;
        RECT 72.680 138.550 72.970 139.625 ;
        RECT 67.905 138.295 68.905 138.325 ;
        RECT 71.435 138.295 72.085 138.325 ;
        RECT 72.675 138.295 72.975 138.550 ;
        RECT 64.705 138.125 66.260 138.190 ;
        RECT 60.310 137.050 60.600 138.125 ;
        RECT 61.195 138.095 62.195 138.125 ;
        RECT 64.725 138.095 65.375 138.125 ;
        RECT 61.595 137.735 61.855 137.780 ;
        RECT 61.195 137.705 62.195 137.735 ;
        RECT 64.725 137.705 65.375 137.735 ;
        RECT 61.175 137.535 65.395 137.705 ;
        RECT 61.195 137.505 62.195 137.535 ;
        RECT 64.725 137.505 65.375 137.535 ;
        RECT 61.595 137.460 61.855 137.505 ;
        RECT 60.760 137.250 60.990 137.395 ;
        RECT 62.400 137.250 62.630 137.395 ;
        RECT 63.330 137.250 63.590 137.325 ;
        RECT 64.335 137.250 64.565 137.395 ;
        RECT 65.535 137.250 65.765 137.395 ;
        RECT 60.760 137.080 65.765 137.250 ;
        RECT 53.595 136.690 55.505 136.795 ;
        RECT 41.065 135.295 42.065 135.325 ;
        RECT 44.595 135.295 45.245 135.325 ;
        RECT 45.835 135.295 46.135 135.550 ;
        RECT 37.865 135.125 39.420 135.190 ;
        RECT 33.470 134.050 33.760 135.125 ;
        RECT 34.355 135.095 35.355 135.125 ;
        RECT 37.885 135.095 38.535 135.125 ;
        RECT 34.335 134.735 34.595 134.780 ;
        RECT 34.335 134.705 35.355 134.735 ;
        RECT 37.885 134.705 38.535 134.735 ;
        RECT 34.335 134.535 38.555 134.705 ;
        RECT 34.335 134.505 35.355 134.535 ;
        RECT 37.885 134.505 38.535 134.535 ;
        RECT 34.335 134.460 34.595 134.505 ;
        RECT 33.920 134.250 34.150 134.395 ;
        RECT 35.560 134.250 35.790 134.395 ;
        RECT 37.495 134.250 37.725 134.395 ;
        RECT 38.295 134.250 38.555 134.325 ;
        RECT 38.695 134.250 38.925 134.395 ;
        RECT 33.920 134.080 38.925 134.250 ;
        RECT 26.755 133.690 28.665 133.795 ;
        RECT 26.760 133.625 28.665 133.690 ;
        RECT 31.155 133.625 32.710 133.795 ;
        RECT 33.465 133.795 33.765 134.050 ;
        RECT 33.920 133.935 34.150 134.080 ;
        RECT 35.560 133.935 35.790 134.080 ;
        RECT 37.495 133.935 37.725 134.080 ;
        RECT 38.295 134.005 38.555 134.080 ;
        RECT 38.695 133.935 38.925 134.080 ;
        RECT 34.355 133.795 35.355 133.825 ;
        RECT 37.885 133.795 38.535 133.825 ;
        RECT 39.130 133.795 39.420 135.125 ;
        RECT 40.180 135.125 42.085 135.295 ;
        RECT 44.575 135.190 46.135 135.295 ;
        RECT 46.890 135.295 47.180 136.625 ;
        RECT 47.775 136.595 48.775 136.625 ;
        RECT 51.305 136.595 51.955 136.625 ;
        RECT 48.595 136.235 48.855 136.280 ;
        RECT 47.775 136.205 48.855 136.235 ;
        RECT 49.910 136.205 50.170 136.280 ;
        RECT 51.305 136.205 51.955 136.235 ;
        RECT 47.755 136.035 51.975 136.205 ;
        RECT 47.775 136.005 48.855 136.035 ;
        RECT 48.595 135.960 48.855 136.005 ;
        RECT 49.910 135.960 50.170 136.035 ;
        RECT 51.305 136.005 51.955 136.035 ;
        RECT 47.340 135.750 47.570 135.895 ;
        RECT 48.980 135.750 49.210 135.895 ;
        RECT 49.880 135.750 50.200 135.795 ;
        RECT 50.915 135.750 51.145 135.895 ;
        RECT 52.115 135.750 52.345 135.895 ;
        RECT 47.340 135.580 52.345 135.750 ;
        RECT 47.340 135.435 47.570 135.580 ;
        RECT 48.980 135.435 49.210 135.580 ;
        RECT 49.880 135.535 50.200 135.580 ;
        RECT 50.915 135.435 51.145 135.580 ;
        RECT 52.115 135.435 52.345 135.580 ;
        RECT 52.550 135.550 52.840 136.625 ;
        RECT 53.600 136.625 55.505 136.690 ;
        RECT 47.775 135.295 48.775 135.325 ;
        RECT 51.305 135.295 51.955 135.325 ;
        RECT 52.545 135.295 52.845 135.550 ;
        RECT 44.575 135.125 46.130 135.190 ;
        RECT 40.180 134.050 40.470 135.125 ;
        RECT 41.065 135.095 42.065 135.125 ;
        RECT 44.595 135.095 45.245 135.125 ;
        RECT 41.065 134.705 42.065 134.735 ;
        RECT 44.595 134.705 45.245 134.735 ;
        RECT 41.045 134.535 45.265 134.705 ;
        RECT 41.065 134.505 42.065 134.535 ;
        RECT 44.595 134.505 45.245 134.535 ;
        RECT 40.630 134.250 40.860 134.395 ;
        RECT 42.270 134.250 42.500 134.395 ;
        RECT 44.205 134.250 44.435 134.395 ;
        RECT 45.405 134.250 45.635 134.395 ;
        RECT 45.840 134.250 46.130 135.125 ;
        RECT 40.630 134.080 46.130 134.250 ;
        RECT 33.465 133.690 35.375 133.795 ;
        RECT 26.760 133.415 27.050 133.625 ;
        RECT 27.645 133.595 28.645 133.625 ;
        RECT 31.175 133.595 31.825 133.625 ;
        RECT 32.420 133.415 32.710 133.625 ;
        RECT 33.470 133.625 35.375 133.690 ;
        RECT 37.865 133.625 39.420 133.795 ;
        RECT 40.175 133.795 40.475 134.050 ;
        RECT 40.630 133.935 40.860 134.080 ;
        RECT 42.270 133.935 42.500 134.080 ;
        RECT 44.205 133.935 44.435 134.080 ;
        RECT 45.405 133.935 45.635 134.080 ;
        RECT 41.065 133.795 42.065 133.825 ;
        RECT 44.595 133.795 45.245 133.825 ;
        RECT 45.840 133.795 46.130 134.080 ;
        RECT 46.890 135.125 48.795 135.295 ;
        RECT 51.285 135.190 52.845 135.295 ;
        RECT 53.600 135.295 53.890 136.625 ;
        RECT 54.485 136.595 55.485 136.625 ;
        RECT 55.730 136.365 55.990 136.685 ;
        RECT 57.995 136.625 59.550 136.795 ;
        RECT 60.305 136.795 60.605 137.050 ;
        RECT 60.760 136.935 60.990 137.080 ;
        RECT 62.400 136.935 62.630 137.080 ;
        RECT 63.330 137.005 63.590 137.080 ;
        RECT 64.335 136.935 64.565 137.080 ;
        RECT 65.535 136.935 65.765 137.080 ;
        RECT 61.195 136.795 62.195 136.825 ;
        RECT 64.725 136.795 65.375 136.825 ;
        RECT 65.970 136.795 66.260 138.125 ;
        RECT 67.020 138.125 68.925 138.295 ;
        RECT 71.415 138.190 72.975 138.295 ;
        RECT 73.730 138.295 74.020 139.690 ;
        RECT 74.595 139.625 75.635 139.795 ;
        RECT 78.125 139.625 79.680 139.795 ;
        RECT 80.435 139.690 80.735 140.050 ;
        RECT 80.890 139.935 81.120 140.080 ;
        RECT 81.725 140.005 81.985 140.080 ;
        RECT 82.530 139.935 82.760 140.080 ;
        RECT 84.465 139.935 84.695 140.080 ;
        RECT 85.665 139.935 85.895 140.080 ;
        RECT 81.325 139.795 82.325 139.825 ;
        RECT 84.855 139.795 85.505 139.825 ;
        RECT 86.100 139.795 86.390 141.125 ;
        RECT 87.150 140.050 87.440 142.625 ;
        RECT 88.035 142.595 89.035 142.625 ;
        RECT 91.565 142.595 92.215 142.625 ;
        RECT 88.035 142.205 89.035 142.235 ;
        RECT 90.170 142.205 90.430 142.280 ;
        RECT 91.565 142.205 92.215 142.235 ;
        RECT 88.015 142.035 92.235 142.205 ;
        RECT 88.035 142.005 89.035 142.035 ;
        RECT 90.170 141.960 90.430 142.035 ;
        RECT 91.565 142.005 92.215 142.035 ;
        RECT 87.600 141.750 87.830 141.895 ;
        RECT 88.015 141.750 88.275 141.825 ;
        RECT 89.240 141.750 89.470 141.895 ;
        RECT 91.175 141.750 91.405 141.895 ;
        RECT 92.375 141.750 92.605 141.895 ;
        RECT 87.600 141.580 92.605 141.750 ;
        RECT 87.600 141.435 87.830 141.580 ;
        RECT 88.015 141.505 88.275 141.580 ;
        RECT 89.240 141.435 89.470 141.580 ;
        RECT 91.175 141.435 91.405 141.580 ;
        RECT 92.375 141.435 92.605 141.580 ;
        RECT 92.810 141.550 93.100 142.625 ;
        RECT 88.035 141.295 89.035 141.325 ;
        RECT 91.565 141.295 92.215 141.325 ;
        RECT 92.805 141.295 93.105 141.550 ;
        RECT 88.015 141.125 89.055 141.295 ;
        RECT 91.545 141.190 93.105 141.295 ;
        RECT 91.545 141.125 93.100 141.190 ;
        RECT 88.035 141.095 89.035 141.125 ;
        RECT 91.565 141.095 92.215 141.125 ;
        RECT 88.450 140.735 88.620 141.095 ;
        RECT 88.035 140.705 89.035 140.735 ;
        RECT 90.170 140.705 90.430 140.780 ;
        RECT 91.565 140.705 92.215 140.735 ;
        RECT 88.015 140.535 89.055 140.705 ;
        RECT 90.170 140.535 92.235 140.705 ;
        RECT 88.035 140.505 89.035 140.535 ;
        RECT 90.170 140.460 90.430 140.535 ;
        RECT 91.565 140.505 92.215 140.535 ;
        RECT 87.600 140.250 87.830 140.395 ;
        RECT 88.435 140.250 88.695 140.325 ;
        RECT 89.240 140.250 89.470 140.395 ;
        RECT 91.175 140.250 91.405 140.395 ;
        RECT 92.375 140.250 92.605 140.395 ;
        RECT 87.600 140.080 92.605 140.250 ;
        RECT 74.615 139.595 75.615 139.625 ;
        RECT 78.145 139.595 78.795 139.625 ;
        RECT 75.030 139.235 75.200 139.595 ;
        RECT 74.615 139.205 75.615 139.235 ;
        RECT 76.750 139.205 77.010 139.280 ;
        RECT 78.145 139.205 78.795 139.235 ;
        RECT 74.595 139.035 75.635 139.205 ;
        RECT 76.750 139.035 78.815 139.205 ;
        RECT 74.615 139.005 75.615 139.035 ;
        RECT 76.750 138.960 77.010 139.035 ;
        RECT 78.145 139.005 78.795 139.035 ;
        RECT 74.180 138.750 74.410 138.895 ;
        RECT 75.820 138.825 76.050 138.895 ;
        RECT 75.820 138.750 76.115 138.825 ;
        RECT 77.755 138.750 77.985 138.895 ;
        RECT 78.955 138.750 79.185 138.895 ;
        RECT 74.180 138.580 79.185 138.750 ;
        RECT 74.180 138.435 74.410 138.580 ;
        RECT 75.820 138.505 76.115 138.580 ;
        RECT 75.820 138.435 76.050 138.505 ;
        RECT 77.755 138.435 77.985 138.580 ;
        RECT 78.955 138.435 79.185 138.580 ;
        RECT 79.390 138.550 79.680 139.625 ;
        RECT 74.615 138.295 75.615 138.325 ;
        RECT 78.145 138.295 78.795 138.325 ;
        RECT 79.385 138.295 79.685 138.550 ;
        RECT 71.415 138.125 72.970 138.190 ;
        RECT 67.020 137.050 67.310 138.125 ;
        RECT 67.905 138.095 68.905 138.125 ;
        RECT 71.435 138.095 72.085 138.125 ;
        RECT 71.845 137.735 72.105 137.780 ;
        RECT 67.905 137.705 68.905 137.735 ;
        RECT 71.435 137.705 72.105 137.735 ;
        RECT 67.885 137.535 72.105 137.705 ;
        RECT 67.905 137.505 68.905 137.535 ;
        RECT 71.435 137.505 72.105 137.535 ;
        RECT 71.845 137.460 72.105 137.505 ;
        RECT 67.470 137.250 67.700 137.395 ;
        RECT 69.110 137.250 69.340 137.395 ;
        RECT 70.040 137.250 70.300 137.325 ;
        RECT 71.045 137.250 71.275 137.395 ;
        RECT 72.245 137.250 72.475 137.395 ;
        RECT 67.470 137.080 72.475 137.250 ;
        RECT 60.305 136.690 62.215 136.795 ;
        RECT 58.015 136.595 58.665 136.625 ;
        RECT 54.485 136.205 55.485 136.235 ;
        RECT 55.775 136.205 55.945 136.365 ;
        RECT 56.620 136.205 56.880 136.280 ;
        RECT 58.015 136.205 58.665 136.235 ;
        RECT 54.465 136.035 58.685 136.205 ;
        RECT 54.485 136.005 55.485 136.035 ;
        RECT 56.620 135.960 56.880 136.035 ;
        RECT 58.015 136.005 58.665 136.035 ;
        RECT 54.050 135.750 54.280 135.895 ;
        RECT 55.690 135.750 55.920 135.895 ;
        RECT 56.590 135.750 56.910 135.795 ;
        RECT 57.625 135.750 57.855 135.895 ;
        RECT 58.825 135.750 59.055 135.895 ;
        RECT 54.050 135.580 59.055 135.750 ;
        RECT 54.050 135.435 54.280 135.580 ;
        RECT 55.690 135.435 55.920 135.580 ;
        RECT 56.590 135.535 56.910 135.580 ;
        RECT 57.625 135.435 57.855 135.580 ;
        RECT 58.825 135.435 59.055 135.580 ;
        RECT 59.260 135.550 59.550 136.625 ;
        RECT 60.310 136.625 62.215 136.690 ;
        RECT 64.705 136.625 66.260 136.795 ;
        RECT 67.015 136.795 67.315 137.050 ;
        RECT 67.470 136.935 67.700 137.080 ;
        RECT 69.110 136.935 69.340 137.080 ;
        RECT 70.040 137.005 70.300 137.080 ;
        RECT 71.045 136.935 71.275 137.080 ;
        RECT 72.245 136.935 72.475 137.080 ;
        RECT 67.905 136.795 68.905 136.825 ;
        RECT 71.435 136.795 72.085 136.825 ;
        RECT 72.680 136.795 72.970 138.125 ;
        RECT 73.730 138.125 75.635 138.295 ;
        RECT 78.125 138.190 79.685 138.295 ;
        RECT 80.440 138.295 80.730 139.690 ;
        RECT 81.305 139.625 82.345 139.795 ;
        RECT 84.835 139.625 86.390 139.795 ;
        RECT 87.145 139.690 87.445 140.050 ;
        RECT 87.600 139.935 87.830 140.080 ;
        RECT 88.435 140.005 88.695 140.080 ;
        RECT 89.240 139.935 89.470 140.080 ;
        RECT 91.175 139.935 91.405 140.080 ;
        RECT 92.375 139.935 92.605 140.080 ;
        RECT 88.035 139.795 89.035 139.825 ;
        RECT 91.565 139.795 92.215 139.825 ;
        RECT 92.810 139.795 93.100 141.125 ;
        RECT 81.325 139.595 82.325 139.625 ;
        RECT 84.855 139.595 85.505 139.625 ;
        RECT 81.740 139.235 81.910 139.595 ;
        RECT 81.325 139.205 82.325 139.235 ;
        RECT 83.460 139.205 83.720 139.280 ;
        RECT 84.855 139.205 85.505 139.235 ;
        RECT 81.305 139.035 82.345 139.205 ;
        RECT 83.460 139.035 85.525 139.205 ;
        RECT 81.325 139.005 82.325 139.035 ;
        RECT 83.460 138.960 83.720 139.035 ;
        RECT 84.855 139.005 85.505 139.035 ;
        RECT 80.890 138.750 81.120 138.895 ;
        RECT 82.530 138.825 82.760 138.895 ;
        RECT 82.530 138.750 82.825 138.825 ;
        RECT 84.465 138.750 84.695 138.895 ;
        RECT 85.665 138.750 85.895 138.895 ;
        RECT 80.890 138.580 85.895 138.750 ;
        RECT 80.890 138.435 81.120 138.580 ;
        RECT 82.530 138.505 82.825 138.580 ;
        RECT 82.530 138.435 82.760 138.505 ;
        RECT 84.465 138.435 84.695 138.580 ;
        RECT 85.665 138.435 85.895 138.580 ;
        RECT 86.100 138.550 86.390 139.625 ;
        RECT 81.325 138.295 82.325 138.325 ;
        RECT 84.855 138.295 85.505 138.325 ;
        RECT 86.095 138.295 86.395 138.550 ;
        RECT 78.125 138.125 79.680 138.190 ;
        RECT 73.730 137.050 74.020 138.125 ;
        RECT 74.615 138.095 75.615 138.125 ;
        RECT 78.145 138.095 78.795 138.125 ;
        RECT 75.015 137.735 75.275 137.780 ;
        RECT 74.615 137.705 75.615 137.735 ;
        RECT 78.145 137.705 78.795 137.735 ;
        RECT 74.595 137.535 78.815 137.705 ;
        RECT 74.615 137.505 75.615 137.535 ;
        RECT 78.145 137.505 78.795 137.535 ;
        RECT 75.015 137.460 75.275 137.505 ;
        RECT 74.180 137.250 74.410 137.395 ;
        RECT 75.820 137.250 76.050 137.395 ;
        RECT 76.750 137.250 77.010 137.325 ;
        RECT 77.755 137.250 77.985 137.395 ;
        RECT 78.955 137.250 79.185 137.395 ;
        RECT 74.180 137.080 79.185 137.250 ;
        RECT 67.015 136.690 68.925 136.795 ;
        RECT 54.485 135.295 55.485 135.325 ;
        RECT 58.015 135.295 58.665 135.325 ;
        RECT 59.255 135.295 59.555 135.550 ;
        RECT 51.285 135.125 52.840 135.190 ;
        RECT 46.890 134.050 47.180 135.125 ;
        RECT 47.775 135.095 48.775 135.125 ;
        RECT 51.305 135.095 51.955 135.125 ;
        RECT 47.755 134.735 48.015 134.780 ;
        RECT 47.755 134.705 48.775 134.735 ;
        RECT 51.305 134.705 51.955 134.735 ;
        RECT 47.755 134.535 51.975 134.705 ;
        RECT 47.755 134.505 48.775 134.535 ;
        RECT 51.305 134.505 51.955 134.535 ;
        RECT 47.755 134.460 48.015 134.505 ;
        RECT 47.340 134.250 47.570 134.395 ;
        RECT 48.980 134.250 49.210 134.395 ;
        RECT 50.915 134.250 51.145 134.395 ;
        RECT 51.715 134.250 51.975 134.325 ;
        RECT 52.115 134.250 52.345 134.395 ;
        RECT 47.340 134.080 52.345 134.250 ;
        RECT 40.175 133.690 42.085 133.795 ;
        RECT 33.470 133.415 33.760 133.625 ;
        RECT 34.355 133.595 35.355 133.625 ;
        RECT 37.885 133.595 38.535 133.625 ;
        RECT 39.130 133.415 39.420 133.625 ;
        RECT 40.180 133.625 42.085 133.690 ;
        RECT 44.575 133.625 46.130 133.795 ;
        RECT 46.885 133.795 47.185 134.050 ;
        RECT 47.340 133.935 47.570 134.080 ;
        RECT 48.980 133.935 49.210 134.080 ;
        RECT 50.915 133.935 51.145 134.080 ;
        RECT 51.715 134.005 51.975 134.080 ;
        RECT 52.115 133.935 52.345 134.080 ;
        RECT 47.775 133.795 48.775 133.825 ;
        RECT 51.305 133.795 51.955 133.825 ;
        RECT 52.550 133.795 52.840 135.125 ;
        RECT 53.600 135.125 55.505 135.295 ;
        RECT 57.995 135.190 59.555 135.295 ;
        RECT 60.310 135.295 60.600 136.625 ;
        RECT 61.195 136.595 62.195 136.625 ;
        RECT 64.725 136.595 65.375 136.625 ;
        RECT 62.015 136.235 62.275 136.280 ;
        RECT 61.195 136.205 62.275 136.235 ;
        RECT 63.330 136.205 63.590 136.280 ;
        RECT 64.725 136.205 65.375 136.235 ;
        RECT 61.175 136.035 65.395 136.205 ;
        RECT 61.195 136.005 62.275 136.035 ;
        RECT 62.015 135.960 62.275 136.005 ;
        RECT 63.330 135.960 63.590 136.035 ;
        RECT 64.725 136.005 65.375 136.035 ;
        RECT 60.760 135.750 60.990 135.895 ;
        RECT 62.400 135.750 62.630 135.895 ;
        RECT 63.300 135.750 63.620 135.795 ;
        RECT 64.335 135.750 64.565 135.895 ;
        RECT 65.535 135.750 65.765 135.895 ;
        RECT 60.760 135.580 65.765 135.750 ;
        RECT 60.760 135.435 60.990 135.580 ;
        RECT 62.400 135.435 62.630 135.580 ;
        RECT 63.300 135.535 63.620 135.580 ;
        RECT 64.335 135.435 64.565 135.580 ;
        RECT 65.535 135.435 65.765 135.580 ;
        RECT 65.970 135.550 66.260 136.625 ;
        RECT 67.020 136.625 68.925 136.690 ;
        RECT 61.195 135.295 62.195 135.325 ;
        RECT 64.725 135.295 65.375 135.325 ;
        RECT 65.965 135.295 66.265 135.550 ;
        RECT 57.995 135.125 59.550 135.190 ;
        RECT 53.600 134.050 53.890 135.125 ;
        RECT 54.485 135.095 55.485 135.125 ;
        RECT 58.015 135.095 58.665 135.125 ;
        RECT 54.485 134.705 55.485 134.735 ;
        RECT 58.015 134.705 58.665 134.735 ;
        RECT 54.465 134.535 58.685 134.705 ;
        RECT 54.485 134.505 55.485 134.535 ;
        RECT 58.015 134.505 58.665 134.535 ;
        RECT 54.050 134.250 54.280 134.395 ;
        RECT 55.690 134.250 55.920 134.395 ;
        RECT 57.625 134.250 57.855 134.395 ;
        RECT 58.825 134.250 59.055 134.395 ;
        RECT 59.260 134.250 59.550 135.125 ;
        RECT 54.050 134.080 59.550 134.250 ;
        RECT 46.885 133.690 48.795 133.795 ;
        RECT 40.180 133.415 40.470 133.625 ;
        RECT 41.065 133.595 42.065 133.625 ;
        RECT 44.595 133.595 45.245 133.625 ;
        RECT 45.840 133.415 46.130 133.625 ;
        RECT 46.890 133.625 48.795 133.690 ;
        RECT 51.285 133.625 52.840 133.795 ;
        RECT 53.595 133.795 53.895 134.050 ;
        RECT 54.050 133.935 54.280 134.080 ;
        RECT 55.690 133.935 55.920 134.080 ;
        RECT 57.625 133.935 57.855 134.080 ;
        RECT 58.825 133.935 59.055 134.080 ;
        RECT 54.485 133.795 55.485 133.825 ;
        RECT 58.015 133.795 58.665 133.825 ;
        RECT 59.260 133.795 59.550 134.080 ;
        RECT 60.310 135.125 62.215 135.295 ;
        RECT 64.705 135.190 66.265 135.295 ;
        RECT 67.020 135.295 67.310 136.625 ;
        RECT 67.905 136.595 68.905 136.625 ;
        RECT 69.150 136.365 69.410 136.685 ;
        RECT 71.415 136.625 72.970 136.795 ;
        RECT 73.725 136.795 74.025 137.050 ;
        RECT 74.180 136.935 74.410 137.080 ;
        RECT 75.820 136.935 76.050 137.080 ;
        RECT 76.750 137.005 77.010 137.080 ;
        RECT 77.755 136.935 77.985 137.080 ;
        RECT 78.955 136.935 79.185 137.080 ;
        RECT 74.615 136.795 75.615 136.825 ;
        RECT 78.145 136.795 78.795 136.825 ;
        RECT 79.390 136.795 79.680 138.125 ;
        RECT 80.440 138.125 82.345 138.295 ;
        RECT 84.835 138.190 86.395 138.295 ;
        RECT 87.150 138.295 87.440 139.690 ;
        RECT 88.015 139.625 89.055 139.795 ;
        RECT 91.545 139.625 93.100 139.795 ;
        RECT 88.035 139.595 89.035 139.625 ;
        RECT 91.565 139.595 92.215 139.625 ;
        RECT 88.450 139.235 88.620 139.595 ;
        RECT 88.035 139.205 89.035 139.235 ;
        RECT 90.170 139.205 90.430 139.280 ;
        RECT 91.565 139.205 92.215 139.235 ;
        RECT 88.015 139.035 89.055 139.205 ;
        RECT 90.170 139.035 92.235 139.205 ;
        RECT 88.035 139.005 89.035 139.035 ;
        RECT 90.170 138.960 90.430 139.035 ;
        RECT 91.565 139.005 92.215 139.035 ;
        RECT 87.600 138.750 87.830 138.895 ;
        RECT 89.240 138.825 89.470 138.895 ;
        RECT 89.240 138.750 89.535 138.825 ;
        RECT 91.175 138.750 91.405 138.895 ;
        RECT 92.375 138.750 92.605 138.895 ;
        RECT 87.600 138.580 92.605 138.750 ;
        RECT 87.600 138.435 87.830 138.580 ;
        RECT 89.240 138.505 89.535 138.580 ;
        RECT 89.240 138.435 89.470 138.505 ;
        RECT 91.175 138.435 91.405 138.580 ;
        RECT 92.375 138.435 92.605 138.580 ;
        RECT 92.810 138.550 93.100 139.625 ;
        RECT 88.035 138.295 89.035 138.325 ;
        RECT 91.565 138.295 92.215 138.325 ;
        RECT 92.805 138.295 93.105 138.550 ;
        RECT 84.835 138.125 86.390 138.190 ;
        RECT 80.440 137.050 80.730 138.125 ;
        RECT 81.325 138.095 82.325 138.125 ;
        RECT 84.855 138.095 85.505 138.125 ;
        RECT 85.265 137.735 85.525 137.780 ;
        RECT 81.325 137.705 82.325 137.735 ;
        RECT 84.855 137.705 85.525 137.735 ;
        RECT 81.305 137.535 85.525 137.705 ;
        RECT 81.325 137.505 82.325 137.535 ;
        RECT 84.855 137.505 85.525 137.535 ;
        RECT 85.265 137.460 85.525 137.505 ;
        RECT 80.890 137.250 81.120 137.395 ;
        RECT 82.530 137.250 82.760 137.395 ;
        RECT 83.460 137.250 83.720 137.325 ;
        RECT 84.465 137.250 84.695 137.395 ;
        RECT 85.665 137.250 85.895 137.395 ;
        RECT 80.890 137.080 85.895 137.250 ;
        RECT 73.725 136.690 75.635 136.795 ;
        RECT 71.435 136.595 72.085 136.625 ;
        RECT 67.905 136.205 68.905 136.235 ;
        RECT 69.195 136.205 69.365 136.365 ;
        RECT 70.040 136.205 70.300 136.280 ;
        RECT 71.435 136.205 72.085 136.235 ;
        RECT 67.885 136.035 72.105 136.205 ;
        RECT 67.905 136.005 68.905 136.035 ;
        RECT 70.040 135.960 70.300 136.035 ;
        RECT 71.435 136.005 72.085 136.035 ;
        RECT 67.470 135.750 67.700 135.895 ;
        RECT 69.110 135.750 69.340 135.895 ;
        RECT 70.010 135.750 70.330 135.795 ;
        RECT 71.045 135.750 71.275 135.895 ;
        RECT 72.245 135.750 72.475 135.895 ;
        RECT 67.470 135.580 72.475 135.750 ;
        RECT 67.470 135.435 67.700 135.580 ;
        RECT 69.110 135.435 69.340 135.580 ;
        RECT 70.010 135.535 70.330 135.580 ;
        RECT 71.045 135.435 71.275 135.580 ;
        RECT 72.245 135.435 72.475 135.580 ;
        RECT 72.680 135.550 72.970 136.625 ;
        RECT 73.730 136.625 75.635 136.690 ;
        RECT 78.125 136.625 79.680 136.795 ;
        RECT 80.435 136.795 80.735 137.050 ;
        RECT 80.890 136.935 81.120 137.080 ;
        RECT 82.530 136.935 82.760 137.080 ;
        RECT 83.460 137.005 83.720 137.080 ;
        RECT 84.465 136.935 84.695 137.080 ;
        RECT 85.665 136.935 85.895 137.080 ;
        RECT 81.325 136.795 82.325 136.825 ;
        RECT 84.855 136.795 85.505 136.825 ;
        RECT 86.100 136.795 86.390 138.125 ;
        RECT 87.150 138.125 89.055 138.295 ;
        RECT 91.545 138.190 93.105 138.295 ;
        RECT 91.545 138.125 93.100 138.190 ;
        RECT 87.150 137.050 87.440 138.125 ;
        RECT 88.035 138.095 89.035 138.125 ;
        RECT 91.565 138.095 92.215 138.125 ;
        RECT 88.435 137.735 88.695 137.780 ;
        RECT 88.035 137.705 89.035 137.735 ;
        RECT 91.565 137.705 92.215 137.735 ;
        RECT 88.015 137.535 92.235 137.705 ;
        RECT 88.035 137.505 89.035 137.535 ;
        RECT 91.565 137.505 92.215 137.535 ;
        RECT 88.435 137.460 88.695 137.505 ;
        RECT 87.600 137.250 87.830 137.395 ;
        RECT 89.240 137.250 89.470 137.395 ;
        RECT 90.170 137.250 90.430 137.325 ;
        RECT 91.175 137.250 91.405 137.395 ;
        RECT 92.375 137.250 92.605 137.395 ;
        RECT 87.600 137.080 92.605 137.250 ;
        RECT 80.435 136.690 82.345 136.795 ;
        RECT 67.905 135.295 68.905 135.325 ;
        RECT 71.435 135.295 72.085 135.325 ;
        RECT 72.675 135.295 72.975 135.550 ;
        RECT 64.705 135.125 66.260 135.190 ;
        RECT 60.310 134.050 60.600 135.125 ;
        RECT 61.195 135.095 62.195 135.125 ;
        RECT 64.725 135.095 65.375 135.125 ;
        RECT 61.175 134.735 61.435 134.780 ;
        RECT 61.175 134.705 62.195 134.735 ;
        RECT 64.725 134.705 65.375 134.735 ;
        RECT 61.175 134.535 65.395 134.705 ;
        RECT 61.175 134.505 62.195 134.535 ;
        RECT 64.725 134.505 65.375 134.535 ;
        RECT 61.175 134.460 61.435 134.505 ;
        RECT 60.760 134.250 60.990 134.395 ;
        RECT 62.400 134.250 62.630 134.395 ;
        RECT 64.335 134.250 64.565 134.395 ;
        RECT 65.135 134.250 65.395 134.325 ;
        RECT 65.535 134.250 65.765 134.395 ;
        RECT 60.760 134.080 65.765 134.250 ;
        RECT 53.595 133.690 55.505 133.795 ;
        RECT 46.890 133.415 47.180 133.625 ;
        RECT 47.775 133.595 48.775 133.625 ;
        RECT 51.305 133.595 51.955 133.625 ;
        RECT 52.550 133.415 52.840 133.625 ;
        RECT 53.600 133.625 55.505 133.690 ;
        RECT 57.995 133.625 59.550 133.795 ;
        RECT 60.305 133.795 60.605 134.050 ;
        RECT 60.760 133.935 60.990 134.080 ;
        RECT 62.400 133.935 62.630 134.080 ;
        RECT 64.335 133.935 64.565 134.080 ;
        RECT 65.135 134.005 65.395 134.080 ;
        RECT 65.535 133.935 65.765 134.080 ;
        RECT 61.195 133.795 62.195 133.825 ;
        RECT 64.725 133.795 65.375 133.825 ;
        RECT 65.970 133.795 66.260 135.125 ;
        RECT 67.020 135.125 68.925 135.295 ;
        RECT 71.415 135.190 72.975 135.295 ;
        RECT 73.730 135.295 74.020 136.625 ;
        RECT 74.615 136.595 75.615 136.625 ;
        RECT 78.145 136.595 78.795 136.625 ;
        RECT 75.435 136.235 75.695 136.280 ;
        RECT 74.615 136.205 75.695 136.235 ;
        RECT 76.750 136.205 77.010 136.280 ;
        RECT 78.145 136.205 78.795 136.235 ;
        RECT 74.595 136.035 78.815 136.205 ;
        RECT 74.615 136.005 75.695 136.035 ;
        RECT 75.435 135.960 75.695 136.005 ;
        RECT 76.750 135.960 77.010 136.035 ;
        RECT 78.145 136.005 78.795 136.035 ;
        RECT 74.180 135.750 74.410 135.895 ;
        RECT 75.820 135.750 76.050 135.895 ;
        RECT 76.720 135.750 77.040 135.795 ;
        RECT 77.755 135.750 77.985 135.895 ;
        RECT 78.955 135.750 79.185 135.895 ;
        RECT 74.180 135.580 79.185 135.750 ;
        RECT 74.180 135.435 74.410 135.580 ;
        RECT 75.820 135.435 76.050 135.580 ;
        RECT 76.720 135.535 77.040 135.580 ;
        RECT 77.755 135.435 77.985 135.580 ;
        RECT 78.955 135.435 79.185 135.580 ;
        RECT 79.390 135.550 79.680 136.625 ;
        RECT 80.440 136.625 82.345 136.690 ;
        RECT 74.615 135.295 75.615 135.325 ;
        RECT 78.145 135.295 78.795 135.325 ;
        RECT 79.385 135.295 79.685 135.550 ;
        RECT 71.415 135.125 72.970 135.190 ;
        RECT 67.020 134.050 67.310 135.125 ;
        RECT 67.905 135.095 68.905 135.125 ;
        RECT 71.435 135.095 72.085 135.125 ;
        RECT 67.905 134.705 68.905 134.735 ;
        RECT 71.435 134.705 72.085 134.735 ;
        RECT 67.885 134.535 72.105 134.705 ;
        RECT 67.905 134.505 68.905 134.535 ;
        RECT 71.435 134.505 72.085 134.535 ;
        RECT 67.470 134.250 67.700 134.395 ;
        RECT 69.110 134.250 69.340 134.395 ;
        RECT 71.045 134.250 71.275 134.395 ;
        RECT 72.245 134.250 72.475 134.395 ;
        RECT 72.680 134.250 72.970 135.125 ;
        RECT 67.470 134.080 72.970 134.250 ;
        RECT 60.305 133.690 62.215 133.795 ;
        RECT 53.600 133.415 53.890 133.625 ;
        RECT 54.485 133.595 55.485 133.625 ;
        RECT 58.015 133.595 58.665 133.625 ;
        RECT 59.260 133.415 59.550 133.625 ;
        RECT 60.310 133.625 62.215 133.690 ;
        RECT 64.705 133.625 66.260 133.795 ;
        RECT 67.015 133.795 67.315 134.050 ;
        RECT 67.470 133.935 67.700 134.080 ;
        RECT 69.110 133.935 69.340 134.080 ;
        RECT 71.045 133.935 71.275 134.080 ;
        RECT 72.245 133.935 72.475 134.080 ;
        RECT 67.905 133.795 68.905 133.825 ;
        RECT 71.435 133.795 72.085 133.825 ;
        RECT 72.680 133.795 72.970 134.080 ;
        RECT 73.730 135.125 75.635 135.295 ;
        RECT 78.125 135.190 79.685 135.295 ;
        RECT 80.440 135.295 80.730 136.625 ;
        RECT 81.325 136.595 82.325 136.625 ;
        RECT 82.570 136.365 82.830 136.685 ;
        RECT 84.835 136.625 86.390 136.795 ;
        RECT 87.145 136.795 87.445 137.050 ;
        RECT 87.600 136.935 87.830 137.080 ;
        RECT 89.240 136.935 89.470 137.080 ;
        RECT 90.170 137.005 90.430 137.080 ;
        RECT 91.175 136.935 91.405 137.080 ;
        RECT 92.375 136.935 92.605 137.080 ;
        RECT 88.035 136.795 89.035 136.825 ;
        RECT 91.565 136.795 92.215 136.825 ;
        RECT 92.810 136.795 93.100 138.125 ;
        RECT 87.145 136.690 89.055 136.795 ;
        RECT 84.855 136.595 85.505 136.625 ;
        RECT 81.325 136.205 82.325 136.235 ;
        RECT 82.615 136.205 82.785 136.365 ;
        RECT 83.460 136.205 83.720 136.280 ;
        RECT 84.855 136.205 85.505 136.235 ;
        RECT 81.305 136.035 85.525 136.205 ;
        RECT 81.325 136.005 82.325 136.035 ;
        RECT 83.460 135.960 83.720 136.035 ;
        RECT 84.855 136.005 85.505 136.035 ;
        RECT 80.890 135.750 81.120 135.895 ;
        RECT 82.530 135.750 82.760 135.895 ;
        RECT 83.430 135.750 83.750 135.795 ;
        RECT 84.465 135.750 84.695 135.895 ;
        RECT 85.665 135.750 85.895 135.895 ;
        RECT 80.890 135.580 85.895 135.750 ;
        RECT 80.890 135.435 81.120 135.580 ;
        RECT 82.530 135.435 82.760 135.580 ;
        RECT 83.430 135.535 83.750 135.580 ;
        RECT 84.465 135.435 84.695 135.580 ;
        RECT 85.665 135.435 85.895 135.580 ;
        RECT 86.100 135.550 86.390 136.625 ;
        RECT 87.150 136.625 89.055 136.690 ;
        RECT 91.545 136.625 93.100 136.795 ;
        RECT 81.325 135.295 82.325 135.325 ;
        RECT 84.855 135.295 85.505 135.325 ;
        RECT 86.095 135.295 86.395 135.550 ;
        RECT 78.125 135.125 79.680 135.190 ;
        RECT 73.730 134.050 74.020 135.125 ;
        RECT 74.615 135.095 75.615 135.125 ;
        RECT 78.145 135.095 78.795 135.125 ;
        RECT 74.595 134.735 74.855 134.780 ;
        RECT 74.595 134.705 75.615 134.735 ;
        RECT 78.145 134.705 78.795 134.735 ;
        RECT 74.595 134.535 78.815 134.705 ;
        RECT 74.595 134.505 75.615 134.535 ;
        RECT 78.145 134.505 78.795 134.535 ;
        RECT 74.595 134.460 74.855 134.505 ;
        RECT 74.180 134.250 74.410 134.395 ;
        RECT 75.820 134.250 76.050 134.395 ;
        RECT 77.755 134.250 77.985 134.395 ;
        RECT 78.555 134.250 78.815 134.325 ;
        RECT 78.955 134.250 79.185 134.395 ;
        RECT 74.180 134.080 79.185 134.250 ;
        RECT 67.015 133.690 68.925 133.795 ;
        RECT 60.310 133.415 60.600 133.625 ;
        RECT 61.195 133.595 62.195 133.625 ;
        RECT 64.725 133.595 65.375 133.625 ;
        RECT 65.970 133.415 66.260 133.625 ;
        RECT 67.020 133.625 68.925 133.690 ;
        RECT 71.415 133.625 72.970 133.795 ;
        RECT 73.725 133.795 74.025 134.050 ;
        RECT 74.180 133.935 74.410 134.080 ;
        RECT 75.820 133.935 76.050 134.080 ;
        RECT 77.755 133.935 77.985 134.080 ;
        RECT 78.555 134.005 78.815 134.080 ;
        RECT 78.955 133.935 79.185 134.080 ;
        RECT 74.615 133.795 75.615 133.825 ;
        RECT 78.145 133.795 78.795 133.825 ;
        RECT 79.390 133.795 79.680 135.125 ;
        RECT 80.440 135.125 82.345 135.295 ;
        RECT 84.835 135.190 86.395 135.295 ;
        RECT 87.150 135.295 87.440 136.625 ;
        RECT 88.035 136.595 89.035 136.625 ;
        RECT 91.565 136.595 92.215 136.625 ;
        RECT 88.855 136.235 89.115 136.280 ;
        RECT 88.035 136.205 89.115 136.235 ;
        RECT 90.170 136.205 90.430 136.280 ;
        RECT 91.565 136.205 92.215 136.235 ;
        RECT 88.015 136.035 92.235 136.205 ;
        RECT 88.035 136.005 89.115 136.035 ;
        RECT 88.855 135.960 89.115 136.005 ;
        RECT 90.170 135.960 90.430 136.035 ;
        RECT 91.565 136.005 92.215 136.035 ;
        RECT 87.600 135.750 87.830 135.895 ;
        RECT 89.240 135.750 89.470 135.895 ;
        RECT 90.140 135.750 90.460 135.795 ;
        RECT 91.175 135.750 91.405 135.895 ;
        RECT 92.375 135.750 92.605 135.895 ;
        RECT 87.600 135.580 92.605 135.750 ;
        RECT 87.600 135.435 87.830 135.580 ;
        RECT 89.240 135.435 89.470 135.580 ;
        RECT 90.140 135.535 90.460 135.580 ;
        RECT 91.175 135.435 91.405 135.580 ;
        RECT 92.375 135.435 92.605 135.580 ;
        RECT 92.810 135.550 93.100 136.625 ;
        RECT 88.035 135.295 89.035 135.325 ;
        RECT 91.565 135.295 92.215 135.325 ;
        RECT 92.805 135.295 93.105 135.550 ;
        RECT 84.835 135.125 86.390 135.190 ;
        RECT 80.440 134.050 80.730 135.125 ;
        RECT 81.325 135.095 82.325 135.125 ;
        RECT 84.855 135.095 85.505 135.125 ;
        RECT 81.325 134.705 82.325 134.735 ;
        RECT 84.855 134.705 85.505 134.735 ;
        RECT 81.305 134.535 85.525 134.705 ;
        RECT 81.325 134.505 82.325 134.535 ;
        RECT 84.855 134.505 85.505 134.535 ;
        RECT 80.890 134.250 81.120 134.395 ;
        RECT 82.530 134.250 82.760 134.395 ;
        RECT 84.465 134.250 84.695 134.395 ;
        RECT 85.665 134.250 85.895 134.395 ;
        RECT 86.100 134.250 86.390 135.125 ;
        RECT 80.890 134.080 86.390 134.250 ;
        RECT 73.725 133.690 75.635 133.795 ;
        RECT 67.020 133.415 67.310 133.625 ;
        RECT 67.905 133.595 68.905 133.625 ;
        RECT 71.435 133.595 72.085 133.625 ;
        RECT 72.680 133.415 72.970 133.625 ;
        RECT 73.730 133.625 75.635 133.690 ;
        RECT 78.125 133.625 79.680 133.795 ;
        RECT 80.435 133.795 80.735 134.050 ;
        RECT 80.890 133.935 81.120 134.080 ;
        RECT 82.530 133.935 82.760 134.080 ;
        RECT 84.465 133.935 84.695 134.080 ;
        RECT 85.665 133.935 85.895 134.080 ;
        RECT 81.325 133.795 82.325 133.825 ;
        RECT 84.855 133.795 85.505 133.825 ;
        RECT 86.100 133.795 86.390 134.080 ;
        RECT 87.150 135.125 89.055 135.295 ;
        RECT 91.545 135.190 93.105 135.295 ;
        RECT 91.545 135.125 93.100 135.190 ;
        RECT 87.150 134.050 87.440 135.125 ;
        RECT 88.035 135.095 89.035 135.125 ;
        RECT 91.565 135.095 92.215 135.125 ;
        RECT 88.015 134.735 88.275 134.780 ;
        RECT 88.015 134.705 89.035 134.735 ;
        RECT 91.565 134.705 92.215 134.735 ;
        RECT 88.015 134.535 92.235 134.705 ;
        RECT 88.015 134.505 89.035 134.535 ;
        RECT 91.565 134.505 92.215 134.535 ;
        RECT 88.015 134.460 88.275 134.505 ;
        RECT 87.600 134.250 87.830 134.395 ;
        RECT 89.240 134.250 89.470 134.395 ;
        RECT 91.175 134.250 91.405 134.395 ;
        RECT 91.975 134.250 92.235 134.325 ;
        RECT 92.375 134.250 92.605 134.395 ;
        RECT 87.600 134.080 92.605 134.250 ;
        RECT 80.435 133.690 82.345 133.795 ;
        RECT 73.730 133.415 74.020 133.625 ;
        RECT 74.615 133.595 75.615 133.625 ;
        RECT 78.145 133.595 78.795 133.625 ;
        RECT 79.390 133.415 79.680 133.625 ;
        RECT 80.440 133.625 82.345 133.690 ;
        RECT 84.835 133.625 86.390 133.795 ;
        RECT 87.145 133.795 87.445 134.050 ;
        RECT 87.600 133.935 87.830 134.080 ;
        RECT 89.240 133.935 89.470 134.080 ;
        RECT 91.175 133.935 91.405 134.080 ;
        RECT 91.975 134.005 92.235 134.080 ;
        RECT 92.375 133.935 92.605 134.080 ;
        RECT 88.035 133.795 89.035 133.825 ;
        RECT 91.565 133.795 92.215 133.825 ;
        RECT 92.810 133.795 93.100 135.125 ;
        RECT 87.145 133.690 89.055 133.795 ;
        RECT 80.440 133.415 80.730 133.625 ;
        RECT 81.325 133.595 82.325 133.625 ;
        RECT 84.855 133.595 85.505 133.625 ;
        RECT 86.100 133.415 86.390 133.625 ;
        RECT 87.150 133.625 89.055 133.690 ;
        RECT 91.545 133.625 93.100 133.795 ;
        RECT 87.150 133.415 87.440 133.625 ;
        RECT 88.035 133.595 89.035 133.625 ;
        RECT 91.565 133.595 92.215 133.625 ;
        RECT 92.810 133.415 93.100 133.625 ;
        RECT 38.295 133.245 38.555 133.320 ;
        RECT 83.040 133.245 83.300 133.320 ;
        RECT 38.295 133.075 83.300 133.245 ;
        RECT 87.210 133.245 87.380 133.415 ;
        RECT 91.975 133.245 92.235 133.320 ;
        RECT 87.210 133.075 92.235 133.245 ;
        RECT 38.295 133.000 38.555 133.075 ;
        RECT 83.040 133.000 83.300 133.075 ;
        RECT 91.975 133.000 92.235 133.075 ;
        RECT 51.715 132.860 51.975 132.935 ;
        RECT 79.975 132.860 80.235 132.935 ;
        RECT 51.715 132.690 80.235 132.860 ;
        RECT 51.715 132.615 51.975 132.690 ;
        RECT 79.975 132.615 80.235 132.690 ;
        RECT 65.135 132.475 65.395 132.550 ;
        RECT 89.750 132.475 90.010 132.550 ;
        RECT 65.135 132.305 90.010 132.475 ;
        RECT 65.135 132.230 65.395 132.305 ;
        RECT 89.750 132.230 90.010 132.305 ;
        RECT 29.780 132.090 30.040 132.165 ;
        RECT 43.200 132.090 43.460 132.165 ;
        RECT 56.590 132.090 56.910 132.135 ;
        RECT 70.040 132.090 70.300 132.165 ;
        RECT 29.780 131.920 70.300 132.090 ;
        RECT 29.780 131.845 30.040 131.920 ;
        RECT 43.200 131.845 43.460 131.920 ;
        RECT 56.590 131.875 56.910 131.920 ;
        RECT 70.040 131.845 70.300 131.920 ;
        RECT 78.555 132.090 78.815 132.165 ;
        RECT 86.685 132.090 86.945 132.165 ;
        RECT 78.555 131.920 86.945 132.090 ;
        RECT 78.555 131.845 78.815 131.920 ;
        RECT 86.685 131.845 86.945 131.920 ;
        RECT 36.490 131.705 36.750 131.780 ;
        RECT 49.910 131.705 50.170 131.780 ;
        RECT 63.330 131.705 63.590 131.780 ;
        RECT 76.750 131.705 77.010 131.780 ;
        RECT 36.490 131.535 77.010 131.705 ;
        RECT 36.490 131.460 36.750 131.535 ;
        RECT 49.910 131.460 50.170 131.535 ;
        RECT 63.330 131.460 63.590 131.535 ;
        RECT 76.750 131.460 77.010 131.535 ;
        RECT 90.125 125.145 90.475 125.175 ;
        RECT 90.125 124.795 108.580 125.145 ;
        RECT 90.125 124.765 90.475 124.795 ;
        RECT 69.995 123.645 70.345 123.675 ;
        RECT 69.995 123.295 110.080 123.645 ;
        RECT 69.995 123.265 70.345 123.295 ;
        RECT 76.705 122.145 77.055 122.175 ;
        RECT 76.705 121.795 111.580 122.145 ;
        RECT 76.705 121.765 77.055 121.795 ;
        RECT 74.350 120.645 74.700 120.675 ;
        RECT 83.415 120.645 83.765 120.675 ;
        RECT 74.350 120.295 113.080 120.645 ;
        RECT 74.350 120.265 74.700 120.295 ;
        RECT 83.415 120.265 83.765 120.295 ;
        RECT 16.010 119.145 16.360 119.175 ;
        RECT 16.010 118.795 114.580 119.145 ;
        RECT 16.010 118.765 16.360 118.795 ;
        RECT 17.510 117.645 17.860 117.675 ;
        RECT 17.510 117.295 116.080 117.645 ;
        RECT 17.510 117.265 17.860 117.295 ;
        RECT 19.010 116.145 19.360 116.175 ;
        RECT 19.010 115.795 117.580 116.145 ;
        RECT 19.010 115.765 19.360 115.795 ;
        RECT 20.510 114.645 20.860 114.675 ;
        RECT 20.510 114.295 119.080 114.645 ;
        RECT 20.510 114.265 20.860 114.295 ;
        RECT 33.745 100.810 34.105 100.815 ;
        RECT 36.745 100.810 37.105 100.815 ;
        RECT 39.745 100.810 40.105 100.815 ;
        RECT 42.745 100.810 43.105 100.815 ;
        RECT 45.745 100.810 46.105 100.815 ;
        RECT 33.470 100.520 46.970 100.810 ;
        RECT 33.680 100.515 34.105 100.520 ;
        RECT 33.680 99.925 33.850 100.515 ;
        RECT 33.990 100.130 34.450 100.360 ;
        RECT 33.650 98.925 33.880 99.925 ;
        RECT 33.680 98.905 33.850 98.925 ;
        RECT 34.135 98.720 34.305 100.130 ;
        RECT 34.590 99.925 34.760 99.945 ;
        RECT 35.180 99.925 35.350 100.520 ;
        RECT 36.680 100.515 37.105 100.520 ;
        RECT 35.490 100.130 35.950 100.360 ;
        RECT 34.560 98.925 34.790 99.925 ;
        RECT 35.150 98.925 35.380 99.925 ;
        RECT 33.990 98.490 34.450 98.720 ;
        RECT 31.900 97.530 32.220 97.790 ;
        RECT 31.515 90.820 31.835 91.080 ;
        RECT 31.590 77.660 31.760 90.820 ;
        RECT 31.975 84.370 32.145 97.530 ;
        RECT 34.135 96.785 34.305 98.490 ;
        RECT 33.990 96.555 34.450 96.785 ;
        RECT 33.680 96.395 33.850 96.415 ;
        RECT 33.650 95.745 33.880 96.395 ;
        RECT 33.680 95.150 33.850 95.745 ;
        RECT 34.135 95.585 34.305 96.555 ;
        RECT 34.590 96.395 34.760 98.925 ;
        RECT 35.180 98.905 35.350 98.925 ;
        RECT 35.635 98.720 35.805 100.130 ;
        RECT 36.090 99.925 36.260 99.945 ;
        RECT 36.680 99.925 36.850 100.515 ;
        RECT 36.990 100.130 37.450 100.360 ;
        RECT 36.060 98.925 36.290 99.925 ;
        RECT 36.650 98.925 36.880 99.925 ;
        RECT 35.490 98.490 35.950 98.720 ;
        RECT 36.090 98.635 36.260 98.925 ;
        RECT 36.680 98.905 36.850 98.925 ;
        RECT 37.135 98.720 37.305 100.130 ;
        RECT 37.590 99.925 37.760 99.945 ;
        RECT 38.180 99.925 38.350 100.520 ;
        RECT 39.745 100.515 40.105 100.520 ;
        RECT 42.680 100.515 43.105 100.520 ;
        RECT 45.745 100.515 46.105 100.520 ;
        RECT 38.490 100.130 38.950 100.360 ;
        RECT 39.990 100.130 40.450 100.360 ;
        RECT 41.490 100.130 41.950 100.360 ;
        RECT 37.560 98.925 37.790 99.925 ;
        RECT 38.150 98.925 38.380 99.925 ;
        RECT 36.420 98.635 36.740 98.680 ;
        RECT 35.635 97.820 35.805 98.490 ;
        RECT 36.090 98.465 36.740 98.635 ;
        RECT 36.990 98.490 37.450 98.720 ;
        RECT 35.590 97.500 35.850 97.820 ;
        RECT 36.090 97.790 36.260 98.465 ;
        RECT 36.420 98.420 36.740 98.465 ;
        RECT 37.135 97.790 37.305 98.490 ;
        RECT 36.015 97.530 36.335 97.790 ;
        RECT 37.060 97.530 37.380 97.790 ;
        RECT 35.635 96.785 35.805 97.500 ;
        RECT 35.490 96.555 35.950 96.785 ;
        RECT 35.180 96.395 35.350 96.415 ;
        RECT 34.560 95.745 34.790 96.395 ;
        RECT 35.150 95.745 35.380 96.395 ;
        RECT 34.590 95.725 34.760 95.745 ;
        RECT 33.990 95.355 34.450 95.585 ;
        RECT 34.135 95.150 34.305 95.355 ;
        RECT 35.180 95.155 35.350 95.745 ;
        RECT 35.635 95.585 35.805 96.555 ;
        RECT 36.090 96.395 36.260 97.530 ;
        RECT 37.135 96.785 37.305 97.530 ;
        RECT 36.990 96.555 37.450 96.785 ;
        RECT 36.680 96.395 36.850 96.415 ;
        RECT 36.060 95.745 36.290 96.395 ;
        RECT 36.650 95.745 36.880 96.395 ;
        RECT 36.090 95.725 36.260 95.745 ;
        RECT 35.490 95.355 35.950 95.585 ;
        RECT 35.180 95.150 35.605 95.155 ;
        RECT 36.680 95.150 36.850 95.745 ;
        RECT 37.135 95.585 37.305 96.555 ;
        RECT 37.590 96.395 37.760 98.925 ;
        RECT 38.180 98.905 38.350 98.925 ;
        RECT 38.635 98.720 38.805 100.130 ;
        RECT 39.090 99.925 39.260 99.945 ;
        RECT 39.680 99.925 39.850 99.945 ;
        RECT 39.060 99.510 39.290 99.925 ;
        RECT 39.650 99.510 39.880 99.925 ;
        RECT 40.135 99.525 40.305 100.130 ;
        RECT 41.635 99.945 41.805 100.130 ;
        RECT 40.590 99.925 40.760 99.945 ;
        RECT 41.180 99.925 41.350 99.945 ;
        RECT 39.060 99.340 39.880 99.510 ;
        RECT 39.060 98.925 39.290 99.340 ;
        RECT 39.650 98.925 39.880 99.340 ;
        RECT 40.060 99.265 40.380 99.525 ;
        RECT 40.560 99.510 40.790 99.925 ;
        RECT 41.150 99.510 41.380 99.925 ;
        RECT 41.560 99.685 41.880 99.945 ;
        RECT 42.090 99.925 42.260 99.945 ;
        RECT 42.680 99.925 42.850 100.515 ;
        RECT 42.990 100.130 43.450 100.360 ;
        RECT 44.490 100.130 44.950 100.360 ;
        RECT 45.990 100.130 46.450 100.360 ;
        RECT 40.560 99.340 41.380 99.510 ;
        RECT 39.090 98.905 39.260 98.925 ;
        RECT 39.680 98.905 39.850 98.925 ;
        RECT 40.135 98.720 40.305 99.265 ;
        RECT 40.560 98.925 40.790 99.340 ;
        RECT 41.150 98.925 41.380 99.340 ;
        RECT 40.590 98.905 40.760 98.925 ;
        RECT 41.180 98.905 41.350 98.925 ;
        RECT 41.635 98.720 41.805 99.685 ;
        RECT 42.060 98.925 42.290 99.925 ;
        RECT 42.650 98.925 42.880 99.925 ;
        RECT 38.490 98.490 38.950 98.720 ;
        RECT 39.990 98.490 40.450 98.720 ;
        RECT 41.490 98.490 41.950 98.720 ;
        RECT 38.560 98.425 38.880 98.490 ;
        RECT 38.635 96.785 38.805 98.425 ;
        RECT 39.015 97.530 39.335 97.790 ;
        RECT 38.490 96.555 38.950 96.785 ;
        RECT 38.180 96.395 38.350 96.415 ;
        RECT 37.560 95.985 37.790 96.395 ;
        RECT 37.515 95.725 37.835 95.985 ;
        RECT 38.150 95.745 38.380 96.395 ;
        RECT 36.990 95.355 37.450 95.585 ;
        RECT 38.180 95.155 38.350 95.745 ;
        RECT 38.635 95.585 38.805 96.555 ;
        RECT 39.090 96.395 39.260 97.530 ;
        RECT 40.135 96.785 40.305 98.490 ;
        RECT 40.515 97.530 40.835 97.790 ;
        RECT 39.990 96.555 40.450 96.785 ;
        RECT 39.680 96.395 39.850 96.415 ;
        RECT 39.060 95.745 39.290 96.395 ;
        RECT 39.650 95.745 39.880 96.395 ;
        RECT 39.090 95.725 39.260 95.745 ;
        RECT 38.490 95.355 38.950 95.585 ;
        RECT 38.180 95.150 38.605 95.155 ;
        RECT 39.680 95.150 39.850 95.745 ;
        RECT 40.135 95.585 40.305 96.555 ;
        RECT 40.590 96.395 40.760 97.530 ;
        RECT 41.635 96.785 41.805 98.490 ;
        RECT 42.090 97.790 42.260 98.925 ;
        RECT 42.680 98.905 42.850 98.925 ;
        RECT 43.135 98.720 43.305 100.130 ;
        RECT 43.590 99.925 43.760 99.945 ;
        RECT 44.180 99.925 44.350 99.945 ;
        RECT 43.560 99.510 43.790 99.925 ;
        RECT 44.150 99.510 44.380 99.925 ;
        RECT 43.560 99.340 44.380 99.510 ;
        RECT 43.560 98.925 43.790 99.340 ;
        RECT 44.150 98.925 44.380 99.340 ;
        RECT 44.635 99.105 44.805 100.130 ;
        RECT 46.135 99.945 46.305 100.130 ;
        RECT 45.090 99.925 45.260 99.945 ;
        RECT 45.680 99.925 45.850 99.945 ;
        RECT 45.060 99.510 45.290 99.925 ;
        RECT 45.650 99.510 45.880 99.925 ;
        RECT 46.060 99.685 46.380 99.945 ;
        RECT 46.590 99.925 46.760 99.945 ;
        RECT 45.060 99.340 45.880 99.510 ;
        RECT 43.590 98.905 43.760 98.925 ;
        RECT 44.180 98.905 44.350 98.925 ;
        RECT 44.560 98.720 44.880 99.105 ;
        RECT 45.060 98.925 45.290 99.340 ;
        RECT 45.650 98.925 45.880 99.340 ;
        RECT 45.090 98.905 45.260 98.925 ;
        RECT 45.680 98.905 45.850 98.925 ;
        RECT 46.135 98.720 46.305 99.685 ;
        RECT 46.560 98.925 46.790 99.925 ;
        RECT 42.990 98.490 43.450 98.720 ;
        RECT 44.490 98.490 44.950 98.720 ;
        RECT 45.990 98.490 46.450 98.720 ;
        RECT 43.060 98.425 43.380 98.490 ;
        RECT 42.015 97.530 42.335 97.790 ;
        RECT 41.490 96.555 41.950 96.785 ;
        RECT 41.180 96.395 41.350 96.415 ;
        RECT 40.560 95.745 40.790 96.395 ;
        RECT 41.150 95.745 41.380 96.395 ;
        RECT 40.590 95.725 40.760 95.745 ;
        RECT 39.990 95.355 40.450 95.585 ;
        RECT 41.180 95.155 41.350 95.745 ;
        RECT 41.635 95.585 41.805 96.555 ;
        RECT 42.090 96.395 42.260 97.530 ;
        RECT 43.135 96.785 43.305 98.425 ;
        RECT 43.515 97.530 43.835 97.790 ;
        RECT 42.990 96.555 43.450 96.785 ;
        RECT 42.680 96.395 42.850 96.415 ;
        RECT 42.060 95.745 42.290 96.395 ;
        RECT 42.650 95.745 42.880 96.395 ;
        RECT 42.090 95.725 42.260 95.745 ;
        RECT 41.490 95.355 41.950 95.585 ;
        RECT 41.180 95.150 41.605 95.155 ;
        RECT 42.680 95.150 42.850 95.745 ;
        RECT 43.135 95.585 43.305 96.555 ;
        RECT 43.590 96.395 43.760 97.530 ;
        RECT 44.635 96.785 44.805 98.490 ;
        RECT 45.015 97.530 45.335 97.790 ;
        RECT 44.490 96.555 44.950 96.785 ;
        RECT 44.180 96.395 44.350 96.415 ;
        RECT 43.560 95.745 43.790 96.395 ;
        RECT 44.150 95.745 44.380 96.395 ;
        RECT 43.590 95.725 43.760 95.745 ;
        RECT 42.990 95.355 43.450 95.585 ;
        RECT 44.180 95.155 44.350 95.745 ;
        RECT 44.635 95.585 44.805 96.555 ;
        RECT 45.090 96.395 45.260 97.530 ;
        RECT 46.135 96.785 46.305 98.490 ;
        RECT 46.590 97.790 46.760 98.925 ;
        RECT 46.515 97.530 46.835 97.790 ;
        RECT 45.990 96.555 46.450 96.785 ;
        RECT 45.680 96.395 45.850 96.415 ;
        RECT 45.060 95.745 45.290 96.395 ;
        RECT 45.650 95.745 45.880 96.395 ;
        RECT 45.090 95.725 45.260 95.745 ;
        RECT 44.490 95.355 44.950 95.585 ;
        RECT 44.180 95.150 44.605 95.155 ;
        RECT 45.680 95.150 45.850 95.745 ;
        RECT 46.135 95.585 46.305 96.555 ;
        RECT 46.590 96.395 46.760 97.530 ;
        RECT 46.560 95.745 46.790 96.395 ;
        RECT 55.445 95.800 69.245 96.090 ;
        RECT 46.590 95.725 46.760 95.745 ;
        RECT 45.990 95.355 46.450 95.585 ;
        RECT 55.905 95.410 56.365 95.640 ;
        RECT 55.535 95.205 55.765 95.210 ;
        RECT 33.470 94.860 46.970 95.150 ;
        RECT 35.245 94.855 35.605 94.860 ;
        RECT 38.245 94.855 38.605 94.860 ;
        RECT 41.245 94.855 41.605 94.860 ;
        RECT 44.245 94.855 44.605 94.860 ;
        RECT 54.480 94.500 55.170 94.530 ;
        RECT 33.470 93.810 55.170 94.500 ;
        RECT 33.680 93.805 34.105 93.810 ;
        RECT 33.680 93.215 33.850 93.805 ;
        RECT 33.990 93.420 34.450 93.650 ;
        RECT 33.650 92.215 33.880 93.215 ;
        RECT 33.680 92.195 33.850 92.215 ;
        RECT 34.135 92.010 34.305 93.420 ;
        RECT 34.515 92.975 34.835 93.235 ;
        RECT 35.180 93.215 35.350 93.810 ;
        RECT 36.680 93.805 37.105 93.810 ;
        RECT 35.490 93.420 35.950 93.650 ;
        RECT 34.560 92.215 34.790 92.975 ;
        RECT 35.150 92.215 35.380 93.215 ;
        RECT 33.990 91.780 34.450 92.010 ;
        RECT 34.135 90.075 34.305 91.780 ;
        RECT 33.990 89.845 34.450 90.075 ;
        RECT 33.680 89.685 33.850 89.705 ;
        RECT 33.055 89.015 33.375 89.275 ;
        RECT 33.650 89.035 33.880 89.685 ;
        RECT 34.135 89.275 34.305 89.845 ;
        RECT 34.590 89.685 34.760 92.215 ;
        RECT 35.180 92.195 35.350 92.215 ;
        RECT 35.635 92.010 35.805 93.420 ;
        RECT 36.090 93.215 36.260 93.235 ;
        RECT 36.680 93.215 36.850 93.805 ;
        RECT 36.990 93.420 37.450 93.650 ;
        RECT 36.060 92.395 36.290 93.215 ;
        RECT 36.015 92.135 36.335 92.395 ;
        RECT 36.650 92.215 36.880 93.215 ;
        RECT 36.680 92.195 36.850 92.215 ;
        RECT 35.490 91.780 35.950 92.010 ;
        RECT 35.635 91.110 35.805 91.780 ;
        RECT 35.590 90.790 35.850 91.110 ;
        RECT 36.090 91.080 36.260 92.135 ;
        RECT 37.135 92.010 37.305 93.420 ;
        RECT 37.590 93.215 37.760 93.235 ;
        RECT 38.180 93.215 38.350 93.810 ;
        RECT 39.745 93.805 40.105 93.810 ;
        RECT 42.680 93.805 43.105 93.810 ;
        RECT 45.745 93.805 46.105 93.810 ;
        RECT 38.490 93.420 38.950 93.650 ;
        RECT 39.990 93.420 40.450 93.650 ;
        RECT 41.490 93.420 41.950 93.650 ;
        RECT 37.560 92.815 37.790 93.215 ;
        RECT 37.515 92.555 37.835 92.815 ;
        RECT 37.560 92.215 37.790 92.555 ;
        RECT 38.150 92.215 38.380 93.215 ;
        RECT 36.990 91.780 37.450 92.010 ;
        RECT 37.135 91.080 37.305 91.780 ;
        RECT 36.015 90.820 36.335 91.080 ;
        RECT 37.060 90.820 37.380 91.080 ;
        RECT 35.635 90.075 35.805 90.790 ;
        RECT 35.490 89.845 35.950 90.075 ;
        RECT 35.180 89.685 35.350 89.705 ;
        RECT 31.900 84.110 32.220 84.370 ;
        RECT 31.515 77.400 31.835 77.660 ;
        RECT 31.590 64.240 31.760 77.400 ;
        RECT 31.975 70.980 32.145 84.110 ;
        RECT 32.670 75.595 32.990 75.855 ;
        RECT 31.930 70.660 32.190 70.980 ;
        RECT 31.515 63.980 31.835 64.240 ;
        RECT 17.510 57.575 17.860 57.605 ;
        RECT 17.510 57.225 28.980 57.575 ;
        RECT 17.510 57.195 17.860 57.225 ;
        RECT 19.010 50.865 19.360 50.895 ;
        RECT 19.010 50.515 28.980 50.865 ;
        RECT 31.590 50.820 31.760 63.980 ;
        RECT 31.975 57.530 32.145 70.660 ;
        RECT 32.285 62.175 32.605 62.435 ;
        RECT 31.900 57.270 32.220 57.530 ;
        RECT 31.515 50.560 31.835 50.820 ;
        RECT 19.010 50.485 19.360 50.515 ;
        RECT 31.900 48.755 32.220 49.015 ;
        RECT 20.510 44.155 20.860 44.185 ;
        RECT 20.510 43.805 28.980 44.155 ;
        RECT 20.510 43.775 20.860 43.805 ;
        RECT 31.975 40.885 32.145 48.755 ;
        RECT 31.900 40.625 32.220 40.885 ;
        RECT 32.360 37.820 32.530 62.175 ;
        RECT 32.745 47.595 32.915 75.595 ;
        RECT 32.670 47.335 32.990 47.595 ;
        RECT 33.130 44.530 33.300 89.015 ;
        RECT 33.680 88.440 33.850 89.035 ;
        RECT 34.060 89.015 34.380 89.275 ;
        RECT 34.560 89.035 34.790 89.685 ;
        RECT 35.150 89.035 35.380 89.685 ;
        RECT 34.590 89.015 34.760 89.035 ;
        RECT 34.135 88.875 34.305 89.015 ;
        RECT 33.990 88.645 34.450 88.875 ;
        RECT 35.180 88.445 35.350 89.035 ;
        RECT 35.635 88.875 35.805 89.845 ;
        RECT 36.090 89.685 36.260 90.820 ;
        RECT 37.135 90.075 37.305 90.820 ;
        RECT 36.990 89.845 37.450 90.075 ;
        RECT 36.680 89.685 36.850 89.705 ;
        RECT 36.060 89.035 36.290 89.685 ;
        RECT 36.650 89.035 36.880 89.685 ;
        RECT 36.090 89.015 36.260 89.035 ;
        RECT 35.490 88.645 35.950 88.875 ;
        RECT 35.180 88.440 35.605 88.445 ;
        RECT 36.680 88.440 36.850 89.035 ;
        RECT 37.135 88.875 37.305 89.845 ;
        RECT 37.590 89.685 37.760 92.215 ;
        RECT 38.180 92.195 38.350 92.215 ;
        RECT 38.635 92.010 38.805 93.420 ;
        RECT 39.090 93.215 39.260 93.235 ;
        RECT 39.680 93.215 39.850 93.235 ;
        RECT 39.060 92.800 39.290 93.215 ;
        RECT 39.650 92.800 39.880 93.215 ;
        RECT 40.135 92.815 40.305 93.420 ;
        RECT 41.635 93.235 41.805 93.420 ;
        RECT 40.590 93.215 40.760 93.235 ;
        RECT 41.180 93.215 41.350 93.235 ;
        RECT 39.060 92.630 39.880 92.800 ;
        RECT 39.060 92.215 39.290 92.630 ;
        RECT 39.650 92.215 39.880 92.630 ;
        RECT 40.060 92.555 40.380 92.815 ;
        RECT 40.560 92.800 40.790 93.215 ;
        RECT 41.150 92.800 41.380 93.215 ;
        RECT 41.560 92.975 41.880 93.235 ;
        RECT 42.090 93.215 42.260 93.235 ;
        RECT 42.680 93.215 42.850 93.805 ;
        RECT 54.480 93.780 55.170 93.810 ;
        RECT 55.535 94.205 55.855 95.205 ;
        RECT 42.990 93.420 43.450 93.650 ;
        RECT 44.490 93.420 44.950 93.650 ;
        RECT 45.990 93.420 46.450 93.650 ;
        RECT 55.535 93.460 55.765 94.205 ;
        RECT 56.020 94.015 56.250 95.410 ;
        RECT 56.505 95.205 56.735 95.800 ;
        RECT 57.285 95.410 57.745 95.640 ;
        RECT 56.415 94.205 56.735 95.205 ;
        RECT 56.915 95.205 57.145 95.210 ;
        RECT 56.915 94.205 57.235 95.205 ;
        RECT 55.905 93.755 56.365 94.015 ;
        RECT 40.560 92.630 41.380 92.800 ;
        RECT 39.090 92.195 39.260 92.215 ;
        RECT 39.680 92.195 39.850 92.215 ;
        RECT 40.135 92.010 40.305 92.555 ;
        RECT 40.560 92.215 40.790 92.630 ;
        RECT 41.150 92.215 41.380 92.630 ;
        RECT 40.590 92.195 40.760 92.215 ;
        RECT 41.180 92.195 41.350 92.215 ;
        RECT 41.635 92.010 41.805 92.975 ;
        RECT 42.060 92.215 42.290 93.215 ;
        RECT 42.650 92.215 42.880 93.215 ;
        RECT 38.490 91.780 38.950 92.010 ;
        RECT 39.990 91.780 40.450 92.010 ;
        RECT 41.490 91.780 41.950 92.010 ;
        RECT 38.560 91.715 38.880 91.780 ;
        RECT 38.635 90.075 38.805 91.715 ;
        RECT 39.015 90.820 39.335 91.080 ;
        RECT 38.490 89.845 38.950 90.075 ;
        RECT 38.180 89.685 38.350 89.705 ;
        RECT 37.560 89.035 37.790 89.685 ;
        RECT 38.150 89.035 38.380 89.685 ;
        RECT 37.590 89.015 37.760 89.035 ;
        RECT 36.990 88.645 37.450 88.875 ;
        RECT 38.180 88.445 38.350 89.035 ;
        RECT 38.635 88.875 38.805 89.845 ;
        RECT 39.090 89.685 39.260 90.820 ;
        RECT 40.135 90.075 40.305 91.780 ;
        RECT 40.515 90.820 40.835 91.080 ;
        RECT 39.990 89.845 40.450 90.075 ;
        RECT 39.680 89.685 39.850 89.705 ;
        RECT 39.060 89.035 39.290 89.685 ;
        RECT 39.650 89.035 39.880 89.685 ;
        RECT 39.090 89.015 39.260 89.035 ;
        RECT 38.490 88.645 38.950 88.875 ;
        RECT 38.180 88.440 38.605 88.445 ;
        RECT 39.680 88.440 39.850 89.035 ;
        RECT 40.135 88.875 40.305 89.845 ;
        RECT 40.590 89.685 40.760 90.820 ;
        RECT 41.635 90.075 41.805 91.780 ;
        RECT 42.090 91.080 42.260 92.215 ;
        RECT 42.680 92.195 42.850 92.215 ;
        RECT 43.135 92.010 43.305 93.420 ;
        RECT 43.590 93.215 43.760 93.235 ;
        RECT 44.180 93.215 44.350 93.235 ;
        RECT 43.560 92.800 43.790 93.215 ;
        RECT 44.150 92.800 44.380 93.215 ;
        RECT 43.560 92.630 44.380 92.800 ;
        RECT 43.560 92.215 43.790 92.630 ;
        RECT 44.150 92.215 44.380 92.630 ;
        RECT 44.635 92.395 44.805 93.420 ;
        RECT 46.135 93.235 46.305 93.420 ;
        RECT 45.090 93.215 45.260 93.235 ;
        RECT 45.680 93.215 45.850 93.235 ;
        RECT 45.060 92.800 45.290 93.215 ;
        RECT 45.650 92.800 45.880 93.215 ;
        RECT 46.060 92.975 46.380 93.235 ;
        RECT 46.590 93.215 46.760 93.235 ;
        RECT 55.535 93.230 56.365 93.460 ;
        RECT 45.060 92.630 45.880 92.800 ;
        RECT 43.590 92.195 43.760 92.215 ;
        RECT 44.180 92.195 44.350 92.215 ;
        RECT 44.560 92.010 44.880 92.395 ;
        RECT 45.060 92.215 45.290 92.630 ;
        RECT 45.650 92.215 45.880 92.630 ;
        RECT 45.090 92.195 45.260 92.215 ;
        RECT 45.680 92.195 45.850 92.215 ;
        RECT 46.135 92.010 46.305 92.975 ;
        RECT 46.560 92.215 46.790 93.215 ;
        RECT 55.535 93.025 55.765 93.030 ;
        RECT 42.990 91.780 43.450 92.010 ;
        RECT 44.490 91.780 44.950 92.010 ;
        RECT 45.990 91.780 46.450 92.010 ;
        RECT 43.060 91.715 43.380 91.780 ;
        RECT 42.015 90.820 42.335 91.080 ;
        RECT 41.490 89.845 41.950 90.075 ;
        RECT 41.180 89.685 41.350 89.705 ;
        RECT 40.560 89.035 40.790 89.685 ;
        RECT 41.150 89.035 41.380 89.685 ;
        RECT 40.590 89.015 40.760 89.035 ;
        RECT 39.990 88.645 40.450 88.875 ;
        RECT 41.180 88.445 41.350 89.035 ;
        RECT 41.635 88.875 41.805 89.845 ;
        RECT 42.090 89.685 42.260 90.820 ;
        RECT 43.135 90.075 43.305 91.715 ;
        RECT 43.515 90.820 43.835 91.080 ;
        RECT 42.990 89.845 43.450 90.075 ;
        RECT 42.680 89.685 42.850 89.705 ;
        RECT 42.060 89.035 42.290 89.685 ;
        RECT 42.650 89.035 42.880 89.685 ;
        RECT 42.090 89.015 42.260 89.035 ;
        RECT 41.490 88.645 41.950 88.875 ;
        RECT 41.180 88.440 41.605 88.445 ;
        RECT 42.680 88.440 42.850 89.035 ;
        RECT 43.135 88.875 43.305 89.845 ;
        RECT 43.590 89.685 43.760 90.820 ;
        RECT 44.635 90.075 44.805 91.780 ;
        RECT 45.015 90.820 45.335 91.080 ;
        RECT 44.490 89.845 44.950 90.075 ;
        RECT 44.180 89.685 44.350 89.705 ;
        RECT 43.560 89.035 43.790 89.685 ;
        RECT 44.150 89.035 44.380 89.685 ;
        RECT 43.590 89.015 43.760 89.035 ;
        RECT 42.990 88.645 43.450 88.875 ;
        RECT 44.180 88.445 44.350 89.035 ;
        RECT 44.635 88.875 44.805 89.845 ;
        RECT 45.090 89.685 45.260 90.820 ;
        RECT 46.135 90.075 46.305 91.780 ;
        RECT 46.590 91.080 46.760 92.215 ;
        RECT 55.535 92.025 55.855 93.025 ;
        RECT 46.515 90.820 46.835 91.080 ;
        RECT 45.990 89.845 46.450 90.075 ;
        RECT 45.680 89.685 45.850 89.705 ;
        RECT 45.060 89.035 45.290 89.685 ;
        RECT 45.650 89.035 45.880 89.685 ;
        RECT 45.090 89.015 45.260 89.035 ;
        RECT 44.490 88.645 44.950 88.875 ;
        RECT 44.180 88.440 44.605 88.445 ;
        RECT 45.680 88.440 45.850 89.035 ;
        RECT 46.135 88.875 46.305 89.845 ;
        RECT 46.590 89.685 46.760 90.820 ;
        RECT 46.560 89.035 46.790 89.685 ;
        RECT 55.535 89.495 55.765 92.025 ;
        RECT 56.020 91.865 56.250 93.230 ;
        RECT 56.505 93.210 56.765 93.530 ;
        RECT 56.915 93.460 57.145 94.205 ;
        RECT 57.400 94.015 57.630 95.410 ;
        RECT 57.885 95.205 58.115 95.800 ;
        RECT 58.665 95.410 59.125 95.640 ;
        RECT 57.795 94.205 58.115 95.205 ;
        RECT 58.295 95.205 58.525 95.210 ;
        RECT 58.295 94.205 58.615 95.205 ;
        RECT 57.285 93.755 57.745 94.015 ;
        RECT 56.915 93.230 57.745 93.460 ;
        RECT 56.505 93.025 56.735 93.210 ;
        RECT 56.415 92.025 56.735 93.025 ;
        RECT 55.905 91.545 56.365 91.865 ;
        RECT 55.905 89.640 56.365 89.900 ;
        RECT 46.590 89.015 46.760 89.035 ;
        RECT 45.990 88.645 46.450 88.875 ;
        RECT 55.535 88.845 55.855 89.495 ;
        RECT 56.020 88.685 56.250 89.640 ;
        RECT 56.505 89.495 56.735 92.025 ;
        RECT 56.415 88.845 56.735 89.495 ;
        RECT 56.915 93.025 57.145 93.030 ;
        RECT 56.915 92.025 57.235 93.025 ;
        RECT 56.915 89.495 57.145 92.025 ;
        RECT 57.400 91.865 57.630 93.230 ;
        RECT 57.885 93.210 58.145 93.530 ;
        RECT 58.295 93.460 58.525 94.205 ;
        RECT 58.780 94.015 59.010 95.410 ;
        RECT 59.265 95.205 59.495 95.800 ;
        RECT 60.045 95.410 60.505 95.640 ;
        RECT 59.175 94.205 59.495 95.205 ;
        RECT 59.675 95.205 59.905 95.210 ;
        RECT 59.675 94.205 59.995 95.205 ;
        RECT 58.665 93.755 59.125 94.015 ;
        RECT 58.295 93.230 59.125 93.460 ;
        RECT 57.885 93.025 58.115 93.210 ;
        RECT 57.795 92.025 58.115 93.025 ;
        RECT 57.285 91.545 57.745 91.865 ;
        RECT 57.285 89.640 57.745 89.900 ;
        RECT 56.915 88.845 57.235 89.495 ;
        RECT 57.400 88.685 57.630 89.640 ;
        RECT 57.885 89.495 58.115 92.025 ;
        RECT 57.795 88.845 58.115 89.495 ;
        RECT 58.295 93.025 58.525 93.030 ;
        RECT 58.295 92.025 58.615 93.025 ;
        RECT 58.295 89.495 58.525 92.025 ;
        RECT 58.780 91.865 59.010 93.230 ;
        RECT 59.265 93.210 59.525 93.530 ;
        RECT 59.675 93.460 59.905 94.205 ;
        RECT 60.160 94.015 60.390 95.410 ;
        RECT 60.645 95.205 60.875 95.800 ;
        RECT 61.425 95.410 61.885 95.640 ;
        RECT 60.555 94.205 60.875 95.205 ;
        RECT 61.055 95.205 61.285 95.210 ;
        RECT 61.055 94.205 61.375 95.205 ;
        RECT 60.045 93.755 60.505 94.015 ;
        RECT 59.675 93.230 60.505 93.460 ;
        RECT 59.265 93.025 59.495 93.210 ;
        RECT 59.175 92.025 59.495 93.025 ;
        RECT 58.665 91.545 59.125 91.865 ;
        RECT 58.665 89.640 59.125 89.900 ;
        RECT 58.295 88.845 58.615 89.495 ;
        RECT 58.780 88.685 59.010 89.640 ;
        RECT 59.265 89.495 59.495 92.025 ;
        RECT 59.175 88.845 59.495 89.495 ;
        RECT 59.675 93.025 59.905 93.030 ;
        RECT 59.675 92.025 59.995 93.025 ;
        RECT 59.675 89.495 59.905 92.025 ;
        RECT 60.160 91.865 60.390 93.230 ;
        RECT 60.645 93.210 60.905 93.530 ;
        RECT 61.055 93.460 61.285 94.205 ;
        RECT 61.540 94.015 61.770 95.410 ;
        RECT 62.025 95.205 62.255 95.800 ;
        RECT 62.805 95.410 63.265 95.640 ;
        RECT 61.935 94.205 62.255 95.205 ;
        RECT 62.435 95.205 62.665 95.210 ;
        RECT 62.435 94.205 62.755 95.205 ;
        RECT 61.425 93.755 61.885 94.015 ;
        RECT 61.055 93.230 61.885 93.460 ;
        RECT 60.645 93.025 60.875 93.210 ;
        RECT 60.555 92.025 60.875 93.025 ;
        RECT 60.045 91.545 60.505 91.865 ;
        RECT 60.045 89.640 60.505 89.900 ;
        RECT 59.675 88.845 59.995 89.495 ;
        RECT 60.160 88.685 60.390 89.640 ;
        RECT 60.645 89.495 60.875 92.025 ;
        RECT 60.555 88.845 60.875 89.495 ;
        RECT 61.055 93.025 61.285 93.030 ;
        RECT 61.055 92.025 61.375 93.025 ;
        RECT 61.055 89.495 61.285 92.025 ;
        RECT 61.540 91.865 61.770 93.230 ;
        RECT 62.025 93.210 62.285 93.530 ;
        RECT 62.435 93.460 62.665 94.205 ;
        RECT 62.920 94.015 63.150 95.410 ;
        RECT 63.405 95.205 63.635 95.800 ;
        RECT 64.185 95.410 64.645 95.640 ;
        RECT 63.315 94.205 63.635 95.205 ;
        RECT 63.815 95.205 64.045 95.210 ;
        RECT 63.815 94.205 64.135 95.205 ;
        RECT 62.805 93.755 63.265 94.015 ;
        RECT 62.435 93.230 63.265 93.460 ;
        RECT 62.025 93.025 62.255 93.210 ;
        RECT 61.935 92.025 62.255 93.025 ;
        RECT 61.425 91.545 61.885 91.865 ;
        RECT 61.425 89.640 61.885 89.900 ;
        RECT 61.055 88.845 61.375 89.495 ;
        RECT 61.540 88.685 61.770 89.640 ;
        RECT 62.025 89.495 62.255 92.025 ;
        RECT 61.935 88.845 62.255 89.495 ;
        RECT 62.435 93.025 62.665 93.030 ;
        RECT 62.435 92.025 62.755 93.025 ;
        RECT 62.435 89.495 62.665 92.025 ;
        RECT 62.920 91.865 63.150 93.230 ;
        RECT 63.405 93.210 63.665 93.530 ;
        RECT 63.815 93.460 64.045 94.205 ;
        RECT 64.300 94.015 64.530 95.410 ;
        RECT 64.785 95.205 65.015 95.800 ;
        RECT 65.565 95.410 66.025 95.640 ;
        RECT 64.695 94.205 65.015 95.205 ;
        RECT 65.195 95.205 65.425 95.210 ;
        RECT 65.195 94.205 65.515 95.205 ;
        RECT 64.185 93.755 64.645 94.015 ;
        RECT 63.815 93.230 64.645 93.460 ;
        RECT 63.405 93.025 63.635 93.210 ;
        RECT 63.315 92.025 63.635 93.025 ;
        RECT 62.805 91.545 63.265 91.865 ;
        RECT 62.805 89.640 63.265 89.900 ;
        RECT 62.435 88.845 62.755 89.495 ;
        RECT 62.920 88.685 63.150 89.640 ;
        RECT 63.405 89.495 63.635 92.025 ;
        RECT 63.315 88.845 63.635 89.495 ;
        RECT 63.815 93.025 64.045 93.030 ;
        RECT 63.815 92.025 64.135 93.025 ;
        RECT 63.815 89.495 64.045 92.025 ;
        RECT 64.300 91.865 64.530 93.230 ;
        RECT 64.785 93.210 65.045 93.530 ;
        RECT 65.195 93.460 65.425 94.205 ;
        RECT 65.680 94.015 65.910 95.410 ;
        RECT 66.165 95.205 66.395 95.800 ;
        RECT 66.945 95.410 67.405 95.640 ;
        RECT 66.075 94.205 66.395 95.205 ;
        RECT 66.575 95.205 66.805 95.210 ;
        RECT 66.575 94.205 66.895 95.205 ;
        RECT 65.565 93.755 66.025 94.015 ;
        RECT 65.195 93.230 66.025 93.460 ;
        RECT 64.785 93.025 65.015 93.210 ;
        RECT 64.695 92.025 65.015 93.025 ;
        RECT 64.185 91.545 64.645 91.865 ;
        RECT 64.185 89.640 64.645 89.900 ;
        RECT 63.815 88.845 64.135 89.495 ;
        RECT 64.300 88.685 64.530 89.640 ;
        RECT 64.785 89.495 65.015 92.025 ;
        RECT 64.695 88.845 65.015 89.495 ;
        RECT 65.195 93.025 65.425 93.030 ;
        RECT 65.195 92.025 65.515 93.025 ;
        RECT 65.195 89.495 65.425 92.025 ;
        RECT 65.680 91.865 65.910 93.230 ;
        RECT 66.165 93.210 66.425 93.530 ;
        RECT 66.575 93.460 66.805 94.205 ;
        RECT 67.060 94.015 67.290 95.410 ;
        RECT 67.545 95.205 67.775 95.800 ;
        RECT 68.325 95.410 68.785 95.640 ;
        RECT 67.455 94.205 67.775 95.205 ;
        RECT 67.955 95.205 68.185 95.210 ;
        RECT 67.955 94.205 68.275 95.205 ;
        RECT 66.945 93.755 67.405 94.015 ;
        RECT 66.575 93.230 67.405 93.460 ;
        RECT 66.165 93.025 66.395 93.210 ;
        RECT 66.075 92.025 66.395 93.025 ;
        RECT 65.565 91.545 66.025 91.865 ;
        RECT 65.565 89.640 66.025 89.900 ;
        RECT 65.195 88.845 65.515 89.495 ;
        RECT 65.680 88.685 65.910 89.640 ;
        RECT 66.165 89.495 66.395 92.025 ;
        RECT 66.075 88.845 66.395 89.495 ;
        RECT 66.575 93.025 66.805 93.030 ;
        RECT 66.575 92.025 66.895 93.025 ;
        RECT 66.575 89.495 66.805 92.025 ;
        RECT 67.060 91.865 67.290 93.230 ;
        RECT 67.545 93.210 67.805 93.530 ;
        RECT 67.955 93.460 68.185 94.205 ;
        RECT 68.440 94.015 68.670 95.410 ;
        RECT 68.925 95.205 69.155 95.800 ;
        RECT 68.835 94.205 69.155 95.205 ;
        RECT 68.325 93.755 68.785 94.015 ;
        RECT 67.955 93.230 68.785 93.460 ;
        RECT 67.545 93.025 67.775 93.210 ;
        RECT 67.455 92.025 67.775 93.025 ;
        RECT 66.945 91.545 67.405 91.865 ;
        RECT 66.945 89.640 67.405 89.900 ;
        RECT 66.575 88.845 66.895 89.495 ;
        RECT 67.060 88.685 67.290 89.640 ;
        RECT 67.545 89.495 67.775 92.025 ;
        RECT 67.455 88.845 67.775 89.495 ;
        RECT 67.955 93.025 68.185 93.030 ;
        RECT 67.955 92.025 68.275 93.025 ;
        RECT 67.955 89.495 68.185 92.025 ;
        RECT 68.440 91.865 68.670 93.230 ;
        RECT 68.925 93.210 69.185 93.530 ;
        RECT 68.925 93.025 69.155 93.210 ;
        RECT 68.835 92.025 69.155 93.025 ;
        RECT 68.325 91.545 68.785 91.865 ;
        RECT 68.325 89.640 68.785 89.900 ;
        RECT 67.955 88.845 68.275 89.495 ;
        RECT 68.440 88.685 68.670 89.640 ;
        RECT 68.925 89.495 69.155 92.025 ;
        RECT 68.835 88.845 69.155 89.495 ;
        RECT 54.480 88.440 55.170 88.470 ;
        RECT 55.905 88.455 56.365 88.685 ;
        RECT 57.285 88.455 57.745 88.685 ;
        RECT 58.665 88.455 59.125 88.685 ;
        RECT 60.045 88.455 60.505 88.685 ;
        RECT 61.425 88.455 61.885 88.685 ;
        RECT 62.805 88.455 63.265 88.685 ;
        RECT 64.185 88.455 64.645 88.685 ;
        RECT 65.565 88.455 66.025 88.685 ;
        RECT 66.945 88.455 67.405 88.685 ;
        RECT 68.325 88.455 68.785 88.685 ;
        RECT 33.470 87.750 55.170 88.440 ;
        RECT 56.020 88.145 56.365 88.455 ;
        RECT 57.400 88.145 57.745 88.455 ;
        RECT 58.780 88.145 59.125 88.455 ;
        RECT 60.160 88.145 60.505 88.455 ;
        RECT 61.540 88.145 61.885 88.455 ;
        RECT 62.920 88.145 63.265 88.455 ;
        RECT 64.300 88.145 64.645 88.455 ;
        RECT 65.680 88.145 66.025 88.455 ;
        RECT 67.060 88.145 67.405 88.455 ;
        RECT 68.440 88.145 68.785 88.455 ;
        RECT 55.905 87.915 56.365 88.145 ;
        RECT 57.285 87.915 57.745 88.145 ;
        RECT 58.665 87.915 59.125 88.145 ;
        RECT 60.045 87.915 60.505 88.145 ;
        RECT 61.425 87.915 61.885 88.145 ;
        RECT 62.805 87.915 63.265 88.145 ;
        RECT 64.185 87.915 64.645 88.145 ;
        RECT 65.565 87.915 66.025 88.145 ;
        RECT 66.945 87.915 67.405 88.145 ;
        RECT 68.325 87.915 68.785 88.145 ;
        RECT 54.480 87.720 55.170 87.750 ;
        RECT 33.745 87.390 34.105 87.395 ;
        RECT 36.745 87.390 37.105 87.395 ;
        RECT 39.745 87.390 40.105 87.395 ;
        RECT 42.745 87.390 43.105 87.395 ;
        RECT 45.745 87.390 46.105 87.395 ;
        RECT 33.470 87.100 46.970 87.390 ;
        RECT 55.535 87.105 55.855 87.755 ;
        RECT 33.680 87.095 34.105 87.100 ;
        RECT 33.680 86.505 33.850 87.095 ;
        RECT 33.990 86.710 34.450 86.940 ;
        RECT 33.650 85.505 33.880 86.505 ;
        RECT 33.680 85.485 33.850 85.505 ;
        RECT 34.135 85.300 34.305 86.710 ;
        RECT 34.590 86.505 34.760 86.525 ;
        RECT 35.180 86.505 35.350 87.100 ;
        RECT 36.680 87.095 37.105 87.100 ;
        RECT 35.490 86.710 35.950 86.940 ;
        RECT 34.560 85.505 34.790 86.505 ;
        RECT 35.150 85.505 35.380 86.505 ;
        RECT 33.990 85.070 34.450 85.300 ;
        RECT 34.135 83.365 34.305 85.070 ;
        RECT 33.990 83.135 34.450 83.365 ;
        RECT 33.680 82.975 33.850 82.995 ;
        RECT 33.650 82.325 33.880 82.975 ;
        RECT 33.680 81.730 33.850 82.325 ;
        RECT 34.135 82.165 34.305 83.135 ;
        RECT 34.590 82.975 34.760 85.505 ;
        RECT 35.180 85.485 35.350 85.505 ;
        RECT 35.635 85.300 35.805 86.710 ;
        RECT 36.090 86.505 36.260 86.525 ;
        RECT 36.680 86.505 36.850 87.095 ;
        RECT 36.990 86.710 37.450 86.940 ;
        RECT 36.060 85.505 36.290 86.505 ;
        RECT 36.650 85.505 36.880 86.505 ;
        RECT 35.490 85.070 35.950 85.300 ;
        RECT 36.090 85.215 36.260 85.505 ;
        RECT 36.680 85.485 36.850 85.505 ;
        RECT 37.135 85.300 37.305 86.710 ;
        RECT 37.590 86.505 37.760 86.525 ;
        RECT 38.180 86.505 38.350 87.100 ;
        RECT 39.745 87.095 40.105 87.100 ;
        RECT 42.680 87.095 43.105 87.100 ;
        RECT 45.745 87.095 46.105 87.100 ;
        RECT 38.490 86.710 38.950 86.940 ;
        RECT 39.990 86.710 40.450 86.940 ;
        RECT 41.490 86.710 41.950 86.940 ;
        RECT 37.560 85.505 37.790 86.505 ;
        RECT 38.150 85.505 38.380 86.505 ;
        RECT 36.420 85.215 36.740 85.260 ;
        RECT 35.635 84.400 35.805 85.070 ;
        RECT 36.090 85.045 36.740 85.215 ;
        RECT 36.990 85.070 37.450 85.300 ;
        RECT 35.590 84.080 35.850 84.400 ;
        RECT 36.090 84.370 36.260 85.045 ;
        RECT 36.420 85.000 36.740 85.045 ;
        RECT 37.135 84.370 37.305 85.070 ;
        RECT 36.015 84.110 36.335 84.370 ;
        RECT 37.060 84.110 37.380 84.370 ;
        RECT 35.635 83.365 35.805 84.080 ;
        RECT 35.490 83.135 35.950 83.365 ;
        RECT 35.180 82.975 35.350 82.995 ;
        RECT 34.560 82.325 34.790 82.975 ;
        RECT 35.150 82.325 35.380 82.975 ;
        RECT 34.590 82.305 34.760 82.325 ;
        RECT 33.990 81.935 34.450 82.165 ;
        RECT 34.135 81.730 34.305 81.935 ;
        RECT 35.180 81.735 35.350 82.325 ;
        RECT 35.635 82.165 35.805 83.135 ;
        RECT 36.090 82.975 36.260 84.110 ;
        RECT 37.135 83.365 37.305 84.110 ;
        RECT 36.990 83.135 37.450 83.365 ;
        RECT 36.680 82.975 36.850 82.995 ;
        RECT 36.060 82.325 36.290 82.975 ;
        RECT 36.650 82.325 36.880 82.975 ;
        RECT 36.090 82.305 36.260 82.325 ;
        RECT 35.490 81.935 35.950 82.165 ;
        RECT 35.180 81.730 35.605 81.735 ;
        RECT 36.680 81.730 36.850 82.325 ;
        RECT 37.135 82.165 37.305 83.135 ;
        RECT 37.590 82.975 37.760 85.505 ;
        RECT 38.180 85.485 38.350 85.505 ;
        RECT 38.635 85.300 38.805 86.710 ;
        RECT 39.090 86.505 39.260 86.525 ;
        RECT 39.680 86.505 39.850 86.525 ;
        RECT 39.060 86.090 39.290 86.505 ;
        RECT 39.650 86.090 39.880 86.505 ;
        RECT 40.135 86.105 40.305 86.710 ;
        RECT 41.635 86.525 41.805 86.710 ;
        RECT 40.590 86.505 40.760 86.525 ;
        RECT 41.180 86.505 41.350 86.525 ;
        RECT 39.060 85.920 39.880 86.090 ;
        RECT 39.060 85.505 39.290 85.920 ;
        RECT 39.650 85.505 39.880 85.920 ;
        RECT 40.060 85.845 40.380 86.105 ;
        RECT 40.560 86.090 40.790 86.505 ;
        RECT 41.150 86.090 41.380 86.505 ;
        RECT 41.560 86.265 41.880 86.525 ;
        RECT 42.090 86.505 42.260 86.525 ;
        RECT 42.680 86.505 42.850 87.095 ;
        RECT 56.020 86.945 56.250 87.915 ;
        RECT 56.415 87.105 56.735 87.755 ;
        RECT 56.915 87.105 57.235 87.755 ;
        RECT 42.990 86.710 43.450 86.940 ;
        RECT 44.490 86.710 44.950 86.940 ;
        RECT 45.990 86.710 46.450 86.940 ;
        RECT 55.905 86.715 56.365 86.945 ;
        RECT 40.560 85.920 41.380 86.090 ;
        RECT 39.090 85.485 39.260 85.505 ;
        RECT 39.680 85.485 39.850 85.505 ;
        RECT 40.135 85.300 40.305 85.845 ;
        RECT 40.560 85.505 40.790 85.920 ;
        RECT 41.150 85.505 41.380 85.920 ;
        RECT 40.590 85.485 40.760 85.505 ;
        RECT 41.180 85.485 41.350 85.505 ;
        RECT 41.635 85.300 41.805 86.265 ;
        RECT 42.060 85.505 42.290 86.505 ;
        RECT 42.650 85.505 42.880 86.505 ;
        RECT 38.490 85.070 38.950 85.300 ;
        RECT 39.990 85.070 40.450 85.300 ;
        RECT 41.490 85.070 41.950 85.300 ;
        RECT 38.560 85.005 38.880 85.070 ;
        RECT 38.635 83.365 38.805 85.005 ;
        RECT 39.015 84.110 39.335 84.370 ;
        RECT 38.490 83.135 38.950 83.365 ;
        RECT 38.180 82.975 38.350 82.995 ;
        RECT 37.560 82.565 37.790 82.975 ;
        RECT 37.515 82.305 37.835 82.565 ;
        RECT 38.150 82.325 38.380 82.975 ;
        RECT 36.990 81.935 37.450 82.165 ;
        RECT 38.180 81.735 38.350 82.325 ;
        RECT 38.635 82.165 38.805 83.135 ;
        RECT 39.090 82.975 39.260 84.110 ;
        RECT 40.135 83.365 40.305 85.070 ;
        RECT 40.515 84.110 40.835 84.370 ;
        RECT 39.990 83.135 40.450 83.365 ;
        RECT 39.680 82.975 39.850 82.995 ;
        RECT 39.060 82.325 39.290 82.975 ;
        RECT 39.650 82.325 39.880 82.975 ;
        RECT 39.090 82.305 39.260 82.325 ;
        RECT 38.490 81.935 38.950 82.165 ;
        RECT 38.180 81.730 38.605 81.735 ;
        RECT 39.680 81.730 39.850 82.325 ;
        RECT 40.135 82.165 40.305 83.135 ;
        RECT 40.590 82.975 40.760 84.110 ;
        RECT 41.635 83.365 41.805 85.070 ;
        RECT 42.090 84.370 42.260 85.505 ;
        RECT 42.680 85.485 42.850 85.505 ;
        RECT 43.135 85.300 43.305 86.710 ;
        RECT 43.590 86.505 43.760 86.525 ;
        RECT 44.180 86.505 44.350 86.525 ;
        RECT 43.560 86.090 43.790 86.505 ;
        RECT 44.150 86.090 44.380 86.505 ;
        RECT 43.560 85.920 44.380 86.090 ;
        RECT 43.560 85.505 43.790 85.920 ;
        RECT 44.150 85.505 44.380 85.920 ;
        RECT 44.635 85.685 44.805 86.710 ;
        RECT 46.135 86.525 46.305 86.710 ;
        RECT 45.090 86.505 45.260 86.525 ;
        RECT 45.680 86.505 45.850 86.525 ;
        RECT 45.060 86.090 45.290 86.505 ;
        RECT 45.650 86.090 45.880 86.505 ;
        RECT 46.060 86.265 46.380 86.525 ;
        RECT 46.590 86.505 46.760 86.525 ;
        RECT 56.505 86.510 56.735 87.105 ;
        RECT 57.400 86.945 57.630 87.915 ;
        RECT 57.795 87.105 58.115 87.755 ;
        RECT 58.295 87.105 58.615 87.755 ;
        RECT 57.285 86.715 57.745 86.945 ;
        RECT 57.885 86.510 58.115 87.105 ;
        RECT 58.780 86.945 59.010 87.915 ;
        RECT 59.175 87.105 59.495 87.755 ;
        RECT 59.675 87.105 59.995 87.755 ;
        RECT 58.665 86.715 59.125 86.945 ;
        RECT 59.265 86.510 59.495 87.105 ;
        RECT 60.160 86.945 60.390 87.915 ;
        RECT 60.555 87.105 60.875 87.755 ;
        RECT 61.055 87.105 61.375 87.755 ;
        RECT 60.045 86.715 60.505 86.945 ;
        RECT 60.645 86.510 60.875 87.105 ;
        RECT 61.540 86.945 61.770 87.915 ;
        RECT 61.935 87.105 62.255 87.755 ;
        RECT 62.435 87.105 62.755 87.755 ;
        RECT 61.425 86.715 61.885 86.945 ;
        RECT 62.025 86.510 62.255 87.105 ;
        RECT 62.920 86.945 63.150 87.915 ;
        RECT 63.315 87.105 63.635 87.755 ;
        RECT 63.815 87.105 64.135 87.755 ;
        RECT 62.805 86.715 63.265 86.945 ;
        RECT 63.405 86.510 63.635 87.105 ;
        RECT 64.300 86.945 64.530 87.915 ;
        RECT 64.695 87.105 65.015 87.755 ;
        RECT 65.195 87.105 65.515 87.755 ;
        RECT 64.185 86.715 64.645 86.945 ;
        RECT 64.785 86.510 65.015 87.105 ;
        RECT 65.680 86.945 65.910 87.915 ;
        RECT 66.075 87.105 66.395 87.755 ;
        RECT 66.575 87.105 66.895 87.755 ;
        RECT 65.565 86.715 66.025 86.945 ;
        RECT 66.165 86.510 66.395 87.105 ;
        RECT 67.060 86.945 67.290 87.915 ;
        RECT 67.455 87.105 67.775 87.755 ;
        RECT 67.955 87.105 68.275 87.755 ;
        RECT 66.945 86.715 67.405 86.945 ;
        RECT 67.545 86.510 67.775 87.105 ;
        RECT 68.440 86.945 68.670 87.915 ;
        RECT 68.835 87.105 69.155 87.755 ;
        RECT 68.325 86.715 68.785 86.945 ;
        RECT 68.925 86.510 69.155 87.105 ;
        RECT 45.060 85.920 45.880 86.090 ;
        RECT 43.590 85.485 43.760 85.505 ;
        RECT 44.180 85.485 44.350 85.505 ;
        RECT 44.560 85.300 44.880 85.685 ;
        RECT 45.060 85.505 45.290 85.920 ;
        RECT 45.650 85.505 45.880 85.920 ;
        RECT 45.090 85.485 45.260 85.505 ;
        RECT 45.680 85.485 45.850 85.505 ;
        RECT 46.135 85.300 46.305 86.265 ;
        RECT 46.560 85.505 46.790 86.505 ;
        RECT 55.445 86.220 69.245 86.510 ;
        RECT 50.600 85.740 50.900 85.770 ;
        RECT 52.260 85.740 52.560 85.770 ;
        RECT 53.920 85.740 54.220 85.770 ;
        RECT 55.580 85.740 55.880 85.770 ;
        RECT 57.240 85.740 57.540 85.770 ;
        RECT 58.900 85.740 59.200 85.770 ;
        RECT 42.990 85.070 43.450 85.300 ;
        RECT 44.490 85.070 44.950 85.300 ;
        RECT 45.990 85.070 46.450 85.300 ;
        RECT 43.060 85.005 43.380 85.070 ;
        RECT 42.015 84.110 42.335 84.370 ;
        RECT 41.490 83.135 41.950 83.365 ;
        RECT 41.180 82.975 41.350 82.995 ;
        RECT 40.560 82.325 40.790 82.975 ;
        RECT 41.150 82.325 41.380 82.975 ;
        RECT 40.590 82.305 40.760 82.325 ;
        RECT 39.990 81.935 40.450 82.165 ;
        RECT 41.180 81.735 41.350 82.325 ;
        RECT 41.635 82.165 41.805 83.135 ;
        RECT 42.090 82.975 42.260 84.110 ;
        RECT 43.135 83.365 43.305 85.005 ;
        RECT 43.515 84.110 43.835 84.370 ;
        RECT 42.990 83.135 43.450 83.365 ;
        RECT 42.680 82.975 42.850 82.995 ;
        RECT 42.060 82.325 42.290 82.975 ;
        RECT 42.650 82.325 42.880 82.975 ;
        RECT 42.090 82.305 42.260 82.325 ;
        RECT 41.490 81.935 41.950 82.165 ;
        RECT 41.180 81.730 41.605 81.735 ;
        RECT 42.680 81.730 42.850 82.325 ;
        RECT 43.135 82.165 43.305 83.135 ;
        RECT 43.590 82.975 43.760 84.110 ;
        RECT 44.635 83.365 44.805 85.070 ;
        RECT 45.015 84.110 45.335 84.370 ;
        RECT 44.490 83.135 44.950 83.365 ;
        RECT 44.180 82.975 44.350 82.995 ;
        RECT 43.560 82.325 43.790 82.975 ;
        RECT 44.150 82.325 44.380 82.975 ;
        RECT 43.590 82.305 43.760 82.325 ;
        RECT 42.990 81.935 43.450 82.165 ;
        RECT 44.180 81.735 44.350 82.325 ;
        RECT 44.635 82.165 44.805 83.135 ;
        RECT 45.090 82.975 45.260 84.110 ;
        RECT 46.135 83.365 46.305 85.070 ;
        RECT 46.590 84.370 46.760 85.505 ;
        RECT 46.515 84.110 46.835 84.370 ;
        RECT 45.990 83.135 46.450 83.365 ;
        RECT 45.680 82.975 45.850 82.995 ;
        RECT 45.060 82.325 45.290 82.975 ;
        RECT 45.650 82.325 45.880 82.975 ;
        RECT 45.090 82.305 45.260 82.325 ;
        RECT 44.490 81.935 44.950 82.165 ;
        RECT 44.180 81.730 44.605 81.735 ;
        RECT 45.680 81.730 45.850 82.325 ;
        RECT 46.135 82.165 46.305 83.135 ;
        RECT 46.590 82.975 46.760 84.110 ;
        RECT 48.940 83.605 49.190 85.710 ;
        RECT 49.720 83.580 50.900 85.740 ;
        RECT 51.380 83.580 52.560 85.740 ;
        RECT 53.040 83.580 54.220 85.740 ;
        RECT 54.700 83.580 55.880 85.740 ;
        RECT 56.360 83.580 57.540 85.740 ;
        RECT 58.020 83.580 59.200 85.740 ;
        RECT 59.680 83.580 60.860 85.740 ;
        RECT 61.340 83.580 62.520 85.740 ;
        RECT 63.000 83.580 64.180 85.740 ;
        RECT 64.660 83.580 65.840 85.740 ;
        RECT 66.320 83.580 67.500 85.740 ;
        RECT 67.980 83.580 69.160 85.740 ;
        RECT 69.690 83.605 69.940 85.710 ;
        RECT 46.560 82.325 46.790 82.975 ;
        RECT 46.590 82.305 46.760 82.325 ;
        RECT 45.990 81.935 46.450 82.165 ;
        RECT 33.470 81.440 46.970 81.730 ;
        RECT 35.245 81.435 35.605 81.440 ;
        RECT 38.245 81.435 38.605 81.440 ;
        RECT 41.245 81.435 41.605 81.440 ;
        RECT 44.245 81.435 44.605 81.440 ;
        RECT 33.745 80.680 34.105 80.685 ;
        RECT 36.745 80.680 37.105 80.685 ;
        RECT 39.745 80.680 40.105 80.685 ;
        RECT 42.745 80.680 43.105 80.685 ;
        RECT 45.745 80.680 46.105 80.685 ;
        RECT 33.470 80.390 46.970 80.680 ;
        RECT 33.680 80.385 34.105 80.390 ;
        RECT 33.680 79.795 33.850 80.385 ;
        RECT 33.990 80.000 34.450 80.230 ;
        RECT 33.650 78.795 33.880 79.795 ;
        RECT 33.680 78.775 33.850 78.795 ;
        RECT 34.135 78.590 34.305 80.000 ;
        RECT 34.515 79.555 34.835 79.815 ;
        RECT 35.180 79.795 35.350 80.390 ;
        RECT 36.680 80.385 37.105 80.390 ;
        RECT 35.490 80.000 35.950 80.230 ;
        RECT 34.560 78.795 34.790 79.555 ;
        RECT 35.150 78.795 35.380 79.795 ;
        RECT 33.990 78.360 34.450 78.590 ;
        RECT 34.135 76.655 34.305 78.360 ;
        RECT 33.990 76.425 34.450 76.655 ;
        RECT 33.680 76.265 33.850 76.285 ;
        RECT 33.650 75.615 33.880 76.265 ;
        RECT 34.135 75.855 34.305 76.425 ;
        RECT 34.590 76.265 34.760 78.795 ;
        RECT 35.180 78.775 35.350 78.795 ;
        RECT 35.635 78.590 35.805 80.000 ;
        RECT 36.090 79.795 36.260 79.815 ;
        RECT 36.680 79.795 36.850 80.385 ;
        RECT 36.990 80.000 37.450 80.230 ;
        RECT 36.060 78.975 36.290 79.795 ;
        RECT 36.015 78.715 36.335 78.975 ;
        RECT 36.650 78.795 36.880 79.795 ;
        RECT 36.680 78.775 36.850 78.795 ;
        RECT 35.490 78.360 35.950 78.590 ;
        RECT 35.635 77.690 35.805 78.360 ;
        RECT 35.590 77.370 35.850 77.690 ;
        RECT 36.090 77.660 36.260 78.715 ;
        RECT 37.135 78.590 37.305 80.000 ;
        RECT 37.590 79.795 37.760 79.815 ;
        RECT 38.180 79.795 38.350 80.390 ;
        RECT 39.745 80.385 40.105 80.390 ;
        RECT 42.680 80.385 43.105 80.390 ;
        RECT 45.745 80.385 46.105 80.390 ;
        RECT 38.490 80.000 38.950 80.230 ;
        RECT 39.990 80.000 40.450 80.230 ;
        RECT 41.490 80.000 41.950 80.230 ;
        RECT 37.560 79.395 37.790 79.795 ;
        RECT 37.515 79.135 37.835 79.395 ;
        RECT 37.560 78.795 37.790 79.135 ;
        RECT 38.150 78.795 38.380 79.795 ;
        RECT 36.990 78.360 37.450 78.590 ;
        RECT 37.135 77.660 37.305 78.360 ;
        RECT 36.015 77.400 36.335 77.660 ;
        RECT 37.060 77.400 37.380 77.660 ;
        RECT 35.635 76.655 35.805 77.370 ;
        RECT 35.490 76.425 35.950 76.655 ;
        RECT 35.180 76.265 35.350 76.285 ;
        RECT 33.680 75.020 33.850 75.615 ;
        RECT 34.060 75.595 34.380 75.855 ;
        RECT 34.560 75.615 34.790 76.265 ;
        RECT 35.150 75.615 35.380 76.265 ;
        RECT 34.590 75.595 34.760 75.615 ;
        RECT 34.135 75.455 34.305 75.595 ;
        RECT 33.990 75.225 34.450 75.455 ;
        RECT 35.180 75.025 35.350 75.615 ;
        RECT 35.635 75.455 35.805 76.425 ;
        RECT 36.090 76.265 36.260 77.400 ;
        RECT 37.135 76.655 37.305 77.400 ;
        RECT 36.990 76.425 37.450 76.655 ;
        RECT 36.680 76.265 36.850 76.285 ;
        RECT 36.060 75.615 36.290 76.265 ;
        RECT 36.650 75.615 36.880 76.265 ;
        RECT 36.090 75.595 36.260 75.615 ;
        RECT 35.490 75.225 35.950 75.455 ;
        RECT 35.180 75.020 35.605 75.025 ;
        RECT 36.680 75.020 36.850 75.615 ;
        RECT 37.135 75.455 37.305 76.425 ;
        RECT 37.590 76.265 37.760 78.795 ;
        RECT 38.180 78.775 38.350 78.795 ;
        RECT 38.635 78.590 38.805 80.000 ;
        RECT 39.090 79.795 39.260 79.815 ;
        RECT 39.680 79.795 39.850 79.815 ;
        RECT 39.060 79.380 39.290 79.795 ;
        RECT 39.650 79.380 39.880 79.795 ;
        RECT 40.135 79.395 40.305 80.000 ;
        RECT 41.635 79.815 41.805 80.000 ;
        RECT 40.590 79.795 40.760 79.815 ;
        RECT 41.180 79.795 41.350 79.815 ;
        RECT 39.060 79.210 39.880 79.380 ;
        RECT 39.060 78.795 39.290 79.210 ;
        RECT 39.650 78.795 39.880 79.210 ;
        RECT 40.060 79.135 40.380 79.395 ;
        RECT 40.560 79.380 40.790 79.795 ;
        RECT 41.150 79.380 41.380 79.795 ;
        RECT 41.560 79.555 41.880 79.815 ;
        RECT 42.090 79.795 42.260 79.815 ;
        RECT 42.680 79.795 42.850 80.385 ;
        RECT 42.990 80.000 43.450 80.230 ;
        RECT 44.490 80.000 44.950 80.230 ;
        RECT 45.990 80.000 46.450 80.230 ;
        RECT 40.560 79.210 41.380 79.380 ;
        RECT 39.090 78.775 39.260 78.795 ;
        RECT 39.680 78.775 39.850 78.795 ;
        RECT 40.135 78.590 40.305 79.135 ;
        RECT 40.560 78.795 40.790 79.210 ;
        RECT 41.150 78.795 41.380 79.210 ;
        RECT 40.590 78.775 40.760 78.795 ;
        RECT 41.180 78.775 41.350 78.795 ;
        RECT 41.635 78.590 41.805 79.555 ;
        RECT 42.060 78.795 42.290 79.795 ;
        RECT 42.650 78.795 42.880 79.795 ;
        RECT 38.490 78.360 38.950 78.590 ;
        RECT 39.990 78.360 40.450 78.590 ;
        RECT 41.490 78.360 41.950 78.590 ;
        RECT 38.560 78.295 38.880 78.360 ;
        RECT 38.635 76.655 38.805 78.295 ;
        RECT 39.015 77.400 39.335 77.660 ;
        RECT 38.490 76.425 38.950 76.655 ;
        RECT 38.180 76.265 38.350 76.285 ;
        RECT 37.560 75.615 37.790 76.265 ;
        RECT 38.150 75.615 38.380 76.265 ;
        RECT 37.590 75.595 37.760 75.615 ;
        RECT 36.990 75.225 37.450 75.455 ;
        RECT 38.180 75.025 38.350 75.615 ;
        RECT 38.635 75.455 38.805 76.425 ;
        RECT 39.090 76.265 39.260 77.400 ;
        RECT 40.135 76.655 40.305 78.360 ;
        RECT 40.515 77.400 40.835 77.660 ;
        RECT 39.990 76.425 40.450 76.655 ;
        RECT 39.680 76.265 39.850 76.285 ;
        RECT 39.060 75.615 39.290 76.265 ;
        RECT 39.650 75.615 39.880 76.265 ;
        RECT 39.090 75.595 39.260 75.615 ;
        RECT 38.490 75.225 38.950 75.455 ;
        RECT 38.180 75.020 38.605 75.025 ;
        RECT 39.680 75.020 39.850 75.615 ;
        RECT 40.135 75.455 40.305 76.425 ;
        RECT 40.590 76.265 40.760 77.400 ;
        RECT 41.635 76.655 41.805 78.360 ;
        RECT 42.090 77.660 42.260 78.795 ;
        RECT 42.680 78.775 42.850 78.795 ;
        RECT 43.135 78.590 43.305 80.000 ;
        RECT 43.590 79.795 43.760 79.815 ;
        RECT 44.180 79.795 44.350 79.815 ;
        RECT 43.560 79.380 43.790 79.795 ;
        RECT 44.150 79.380 44.380 79.795 ;
        RECT 43.560 79.210 44.380 79.380 ;
        RECT 43.560 78.795 43.790 79.210 ;
        RECT 44.150 78.795 44.380 79.210 ;
        RECT 44.635 78.975 44.805 80.000 ;
        RECT 46.135 79.815 46.305 80.000 ;
        RECT 45.090 79.795 45.260 79.815 ;
        RECT 45.680 79.795 45.850 79.815 ;
        RECT 45.060 79.380 45.290 79.795 ;
        RECT 45.650 79.380 45.880 79.795 ;
        RECT 46.060 79.555 46.380 79.815 ;
        RECT 46.590 79.795 46.760 79.815 ;
        RECT 45.060 79.210 45.880 79.380 ;
        RECT 43.590 78.775 43.760 78.795 ;
        RECT 44.180 78.775 44.350 78.795 ;
        RECT 44.560 78.590 44.880 78.975 ;
        RECT 45.060 78.795 45.290 79.210 ;
        RECT 45.650 78.795 45.880 79.210 ;
        RECT 45.090 78.775 45.260 78.795 ;
        RECT 45.680 78.775 45.850 78.795 ;
        RECT 46.135 78.590 46.305 79.555 ;
        RECT 46.560 78.795 46.790 79.795 ;
        RECT 42.990 78.360 43.450 78.590 ;
        RECT 44.490 78.360 44.950 78.590 ;
        RECT 45.990 78.360 46.450 78.590 ;
        RECT 43.060 78.295 43.380 78.360 ;
        RECT 42.015 77.400 42.335 77.660 ;
        RECT 41.490 76.425 41.950 76.655 ;
        RECT 41.180 76.265 41.350 76.285 ;
        RECT 40.560 75.615 40.790 76.265 ;
        RECT 41.150 75.615 41.380 76.265 ;
        RECT 40.590 75.595 40.760 75.615 ;
        RECT 39.990 75.225 40.450 75.455 ;
        RECT 41.180 75.025 41.350 75.615 ;
        RECT 41.635 75.455 41.805 76.425 ;
        RECT 42.090 76.265 42.260 77.400 ;
        RECT 43.135 76.655 43.305 78.295 ;
        RECT 43.515 77.400 43.835 77.660 ;
        RECT 42.990 76.425 43.450 76.655 ;
        RECT 42.680 76.265 42.850 76.285 ;
        RECT 42.060 75.615 42.290 76.265 ;
        RECT 42.650 75.615 42.880 76.265 ;
        RECT 42.090 75.595 42.260 75.615 ;
        RECT 41.490 75.225 41.950 75.455 ;
        RECT 41.180 75.020 41.605 75.025 ;
        RECT 42.680 75.020 42.850 75.615 ;
        RECT 43.135 75.455 43.305 76.425 ;
        RECT 43.590 76.265 43.760 77.400 ;
        RECT 44.635 76.655 44.805 78.360 ;
        RECT 45.015 77.400 45.335 77.660 ;
        RECT 44.490 76.425 44.950 76.655 ;
        RECT 44.180 76.265 44.350 76.285 ;
        RECT 43.560 75.615 43.790 76.265 ;
        RECT 44.150 75.615 44.380 76.265 ;
        RECT 43.590 75.595 43.760 75.615 ;
        RECT 42.990 75.225 43.450 75.455 ;
        RECT 44.180 75.025 44.350 75.615 ;
        RECT 44.635 75.455 44.805 76.425 ;
        RECT 45.090 76.265 45.260 77.400 ;
        RECT 46.135 76.655 46.305 78.360 ;
        RECT 46.590 77.660 46.760 78.795 ;
        RECT 46.515 77.400 46.835 77.660 ;
        RECT 45.990 76.425 46.450 76.655 ;
        RECT 45.680 76.265 45.850 76.285 ;
        RECT 45.060 75.615 45.290 76.265 ;
        RECT 45.650 75.615 45.880 76.265 ;
        RECT 45.090 75.595 45.260 75.615 ;
        RECT 44.490 75.225 44.950 75.455 ;
        RECT 44.180 75.020 44.605 75.025 ;
        RECT 45.680 75.020 45.850 75.615 ;
        RECT 46.135 75.455 46.305 76.425 ;
        RECT 46.590 76.265 46.760 77.400 ;
        RECT 46.560 75.615 46.790 76.265 ;
        RECT 46.590 75.595 46.760 75.615 ;
        RECT 45.990 75.225 46.450 75.455 ;
        RECT 33.470 74.730 46.970 75.020 ;
        RECT 35.245 74.725 35.605 74.730 ;
        RECT 38.245 74.725 38.605 74.730 ;
        RECT 41.245 74.725 41.605 74.730 ;
        RECT 44.245 74.725 44.605 74.730 ;
        RECT 33.745 73.970 34.105 73.975 ;
        RECT 36.745 73.970 37.105 73.975 ;
        RECT 39.745 73.970 40.105 73.975 ;
        RECT 42.745 73.970 43.105 73.975 ;
        RECT 45.745 73.970 46.105 73.975 ;
        RECT 33.470 73.680 46.970 73.970 ;
        RECT 33.680 73.675 34.105 73.680 ;
        RECT 33.680 73.085 33.850 73.675 ;
        RECT 33.990 73.290 34.450 73.520 ;
        RECT 33.650 72.085 33.880 73.085 ;
        RECT 33.680 72.065 33.850 72.085 ;
        RECT 34.135 71.880 34.305 73.290 ;
        RECT 34.590 73.085 34.760 73.105 ;
        RECT 35.180 73.085 35.350 73.680 ;
        RECT 36.680 73.675 37.105 73.680 ;
        RECT 35.490 73.290 35.950 73.520 ;
        RECT 34.560 72.085 34.790 73.085 ;
        RECT 35.150 72.085 35.380 73.085 ;
        RECT 33.990 71.650 34.450 71.880 ;
        RECT 34.135 69.945 34.305 71.650 ;
        RECT 33.990 69.715 34.450 69.945 ;
        RECT 33.680 69.555 33.850 69.575 ;
        RECT 33.650 68.905 33.880 69.555 ;
        RECT 33.680 68.310 33.850 68.905 ;
        RECT 34.135 68.745 34.305 69.715 ;
        RECT 34.590 69.555 34.760 72.085 ;
        RECT 35.180 72.065 35.350 72.085 ;
        RECT 35.635 71.880 35.805 73.290 ;
        RECT 36.090 73.085 36.260 73.105 ;
        RECT 36.680 73.085 36.850 73.675 ;
        RECT 36.990 73.290 37.450 73.520 ;
        RECT 36.060 72.085 36.290 73.085 ;
        RECT 36.650 72.085 36.880 73.085 ;
        RECT 35.490 71.650 35.950 71.880 ;
        RECT 36.090 71.795 36.260 72.085 ;
        RECT 36.680 72.065 36.850 72.085 ;
        RECT 37.135 71.880 37.305 73.290 ;
        RECT 37.590 73.085 37.760 73.105 ;
        RECT 38.180 73.085 38.350 73.680 ;
        RECT 39.745 73.675 40.105 73.680 ;
        RECT 42.680 73.675 43.105 73.680 ;
        RECT 45.745 73.675 46.105 73.680 ;
        RECT 38.490 73.290 38.950 73.520 ;
        RECT 39.990 73.290 40.450 73.520 ;
        RECT 41.490 73.290 41.950 73.520 ;
        RECT 37.560 72.085 37.790 73.085 ;
        RECT 38.150 72.085 38.380 73.085 ;
        RECT 36.420 71.795 36.740 71.840 ;
        RECT 35.635 70.980 35.805 71.650 ;
        RECT 36.090 71.625 36.740 71.795 ;
        RECT 36.990 71.650 37.450 71.880 ;
        RECT 35.590 70.660 35.850 70.980 ;
        RECT 36.090 70.950 36.260 71.625 ;
        RECT 36.420 71.580 36.740 71.625 ;
        RECT 37.135 70.950 37.305 71.650 ;
        RECT 36.015 70.690 36.335 70.950 ;
        RECT 37.060 70.690 37.380 70.950 ;
        RECT 35.635 69.945 35.805 70.660 ;
        RECT 35.490 69.715 35.950 69.945 ;
        RECT 35.180 69.555 35.350 69.575 ;
        RECT 34.560 68.905 34.790 69.555 ;
        RECT 35.150 68.905 35.380 69.555 ;
        RECT 34.590 68.885 34.760 68.905 ;
        RECT 33.990 68.515 34.450 68.745 ;
        RECT 34.135 68.310 34.305 68.515 ;
        RECT 35.180 68.315 35.350 68.905 ;
        RECT 35.635 68.745 35.805 69.715 ;
        RECT 36.090 69.555 36.260 70.690 ;
        RECT 37.135 69.945 37.305 70.690 ;
        RECT 36.990 69.715 37.450 69.945 ;
        RECT 36.680 69.555 36.850 69.575 ;
        RECT 36.060 68.905 36.290 69.555 ;
        RECT 36.650 68.905 36.880 69.555 ;
        RECT 36.090 68.885 36.260 68.905 ;
        RECT 35.490 68.515 35.950 68.745 ;
        RECT 35.180 68.310 35.605 68.315 ;
        RECT 36.680 68.310 36.850 68.905 ;
        RECT 37.135 68.745 37.305 69.715 ;
        RECT 37.590 69.555 37.760 72.085 ;
        RECT 38.180 72.065 38.350 72.085 ;
        RECT 38.635 71.880 38.805 73.290 ;
        RECT 39.090 73.085 39.260 73.105 ;
        RECT 39.680 73.085 39.850 73.105 ;
        RECT 39.060 72.670 39.290 73.085 ;
        RECT 39.650 72.670 39.880 73.085 ;
        RECT 40.135 72.685 40.305 73.290 ;
        RECT 41.635 73.105 41.805 73.290 ;
        RECT 40.590 73.085 40.760 73.105 ;
        RECT 41.180 73.085 41.350 73.105 ;
        RECT 39.060 72.500 39.880 72.670 ;
        RECT 39.060 72.085 39.290 72.500 ;
        RECT 39.650 72.085 39.880 72.500 ;
        RECT 40.060 72.425 40.380 72.685 ;
        RECT 40.560 72.670 40.790 73.085 ;
        RECT 41.150 72.670 41.380 73.085 ;
        RECT 41.560 72.845 41.880 73.105 ;
        RECT 42.090 73.085 42.260 73.105 ;
        RECT 42.680 73.085 42.850 73.675 ;
        RECT 42.990 73.290 43.450 73.520 ;
        RECT 44.490 73.290 44.950 73.520 ;
        RECT 45.990 73.290 46.450 73.520 ;
        RECT 40.560 72.500 41.380 72.670 ;
        RECT 39.090 72.065 39.260 72.085 ;
        RECT 39.680 72.065 39.850 72.085 ;
        RECT 40.135 71.880 40.305 72.425 ;
        RECT 40.560 72.085 40.790 72.500 ;
        RECT 41.150 72.085 41.380 72.500 ;
        RECT 40.590 72.065 40.760 72.085 ;
        RECT 41.180 72.065 41.350 72.085 ;
        RECT 41.635 71.880 41.805 72.845 ;
        RECT 42.060 72.085 42.290 73.085 ;
        RECT 42.650 72.085 42.880 73.085 ;
        RECT 38.490 71.650 38.950 71.880 ;
        RECT 39.990 71.650 40.450 71.880 ;
        RECT 41.490 71.650 41.950 71.880 ;
        RECT 38.560 71.585 38.880 71.650 ;
        RECT 38.635 69.945 38.805 71.585 ;
        RECT 39.015 70.690 39.335 70.950 ;
        RECT 38.490 69.715 38.950 69.945 ;
        RECT 38.180 69.555 38.350 69.575 ;
        RECT 37.560 69.145 37.790 69.555 ;
        RECT 37.515 68.885 37.835 69.145 ;
        RECT 38.150 68.905 38.380 69.555 ;
        RECT 36.990 68.515 37.450 68.745 ;
        RECT 38.180 68.315 38.350 68.905 ;
        RECT 38.635 68.745 38.805 69.715 ;
        RECT 39.090 69.555 39.260 70.690 ;
        RECT 40.135 69.945 40.305 71.650 ;
        RECT 40.515 70.690 40.835 70.950 ;
        RECT 39.990 69.715 40.450 69.945 ;
        RECT 39.680 69.555 39.850 69.575 ;
        RECT 39.060 68.905 39.290 69.555 ;
        RECT 39.650 68.905 39.880 69.555 ;
        RECT 39.090 68.885 39.260 68.905 ;
        RECT 38.490 68.515 38.950 68.745 ;
        RECT 38.180 68.310 38.605 68.315 ;
        RECT 39.680 68.310 39.850 68.905 ;
        RECT 40.135 68.745 40.305 69.715 ;
        RECT 40.590 69.555 40.760 70.690 ;
        RECT 41.635 69.945 41.805 71.650 ;
        RECT 42.090 70.950 42.260 72.085 ;
        RECT 42.680 72.065 42.850 72.085 ;
        RECT 43.135 71.880 43.305 73.290 ;
        RECT 43.590 73.085 43.760 73.105 ;
        RECT 44.180 73.085 44.350 73.105 ;
        RECT 43.560 72.670 43.790 73.085 ;
        RECT 44.150 72.670 44.380 73.085 ;
        RECT 43.560 72.500 44.380 72.670 ;
        RECT 43.560 72.085 43.790 72.500 ;
        RECT 44.150 72.085 44.380 72.500 ;
        RECT 44.635 72.265 44.805 73.290 ;
        RECT 46.135 73.105 46.305 73.290 ;
        RECT 45.090 73.085 45.260 73.105 ;
        RECT 45.680 73.085 45.850 73.105 ;
        RECT 45.060 72.670 45.290 73.085 ;
        RECT 45.650 72.670 45.880 73.085 ;
        RECT 46.060 72.845 46.380 73.105 ;
        RECT 46.590 73.085 46.760 73.105 ;
        RECT 45.060 72.500 45.880 72.670 ;
        RECT 43.590 72.065 43.760 72.085 ;
        RECT 44.180 72.065 44.350 72.085 ;
        RECT 44.560 71.880 44.880 72.265 ;
        RECT 45.060 72.085 45.290 72.500 ;
        RECT 45.650 72.085 45.880 72.500 ;
        RECT 45.090 72.065 45.260 72.085 ;
        RECT 45.680 72.065 45.850 72.085 ;
        RECT 46.135 71.880 46.305 72.845 ;
        RECT 46.560 72.085 46.790 73.085 ;
        RECT 102.225 72.950 103.405 75.110 ;
        RECT 103.885 72.950 105.065 75.110 ;
        RECT 105.545 72.950 106.725 75.110 ;
        RECT 107.205 72.950 108.385 75.110 ;
        RECT 108.865 72.950 110.045 75.110 ;
        RECT 110.525 72.950 111.705 75.110 ;
        RECT 112.185 72.950 113.365 75.110 ;
        RECT 113.845 72.950 115.025 75.110 ;
        RECT 115.505 72.950 116.685 75.110 ;
        RECT 117.165 72.950 118.345 75.110 ;
        RECT 118.825 72.950 120.005 75.110 ;
        RECT 120.485 72.950 121.665 75.110 ;
        RECT 42.990 71.650 43.450 71.880 ;
        RECT 44.490 71.650 44.950 71.880 ;
        RECT 45.990 71.650 46.450 71.880 ;
        RECT 43.060 71.585 43.380 71.650 ;
        RECT 42.015 70.690 42.335 70.950 ;
        RECT 41.490 69.715 41.950 69.945 ;
        RECT 41.180 69.555 41.350 69.575 ;
        RECT 40.560 68.905 40.790 69.555 ;
        RECT 41.150 68.905 41.380 69.555 ;
        RECT 40.590 68.885 40.760 68.905 ;
        RECT 39.990 68.515 40.450 68.745 ;
        RECT 41.180 68.315 41.350 68.905 ;
        RECT 41.635 68.745 41.805 69.715 ;
        RECT 42.090 69.555 42.260 70.690 ;
        RECT 43.135 69.945 43.305 71.585 ;
        RECT 43.515 70.690 43.835 70.950 ;
        RECT 42.990 69.715 43.450 69.945 ;
        RECT 42.680 69.555 42.850 69.575 ;
        RECT 42.060 68.905 42.290 69.555 ;
        RECT 42.650 68.905 42.880 69.555 ;
        RECT 42.090 68.885 42.260 68.905 ;
        RECT 41.490 68.515 41.950 68.745 ;
        RECT 41.180 68.310 41.605 68.315 ;
        RECT 42.680 68.310 42.850 68.905 ;
        RECT 43.135 68.745 43.305 69.715 ;
        RECT 43.590 69.555 43.760 70.690 ;
        RECT 44.635 69.945 44.805 71.650 ;
        RECT 45.015 70.690 45.335 70.950 ;
        RECT 44.490 69.715 44.950 69.945 ;
        RECT 44.180 69.555 44.350 69.575 ;
        RECT 43.560 68.905 43.790 69.555 ;
        RECT 44.150 68.905 44.380 69.555 ;
        RECT 43.590 68.885 43.760 68.905 ;
        RECT 42.990 68.515 43.450 68.745 ;
        RECT 44.180 68.315 44.350 68.905 ;
        RECT 44.635 68.745 44.805 69.715 ;
        RECT 45.090 69.555 45.260 70.690 ;
        RECT 46.135 69.945 46.305 71.650 ;
        RECT 46.590 70.950 46.760 72.085 ;
        RECT 46.515 70.690 46.835 70.950 ;
        RECT 45.990 69.715 46.450 69.945 ;
        RECT 45.680 69.555 45.850 69.575 ;
        RECT 45.060 68.905 45.290 69.555 ;
        RECT 45.650 68.905 45.880 69.555 ;
        RECT 45.090 68.885 45.260 68.905 ;
        RECT 44.490 68.515 44.950 68.745 ;
        RECT 44.180 68.310 44.605 68.315 ;
        RECT 45.680 68.310 45.850 68.905 ;
        RECT 46.135 68.745 46.305 69.715 ;
        RECT 46.590 69.555 46.760 70.690 ;
        RECT 46.560 68.905 46.790 69.555 ;
        RECT 46.590 68.885 46.760 68.905 ;
        RECT 45.990 68.515 46.450 68.745 ;
        RECT 33.470 68.020 46.970 68.310 ;
        RECT 35.245 68.015 35.605 68.020 ;
        RECT 38.245 68.015 38.605 68.020 ;
        RECT 41.245 68.015 41.605 68.020 ;
        RECT 44.245 68.015 44.605 68.020 ;
        RECT 33.745 67.260 34.105 67.265 ;
        RECT 36.745 67.260 37.105 67.265 ;
        RECT 39.745 67.260 40.105 67.265 ;
        RECT 42.745 67.260 43.105 67.265 ;
        RECT 45.745 67.260 46.105 67.265 ;
        RECT 33.470 66.970 46.970 67.260 ;
        RECT 33.680 66.965 34.105 66.970 ;
        RECT 33.680 66.375 33.850 66.965 ;
        RECT 33.990 66.580 34.450 66.810 ;
        RECT 33.650 65.375 33.880 66.375 ;
        RECT 33.680 65.355 33.850 65.375 ;
        RECT 34.135 65.170 34.305 66.580 ;
        RECT 34.515 66.135 34.835 66.395 ;
        RECT 35.180 66.375 35.350 66.970 ;
        RECT 36.680 66.965 37.105 66.970 ;
        RECT 35.490 66.580 35.950 66.810 ;
        RECT 34.560 65.375 34.790 66.135 ;
        RECT 35.150 65.375 35.380 66.375 ;
        RECT 33.990 64.940 34.450 65.170 ;
        RECT 34.135 63.235 34.305 64.940 ;
        RECT 33.990 63.005 34.450 63.235 ;
        RECT 33.680 62.845 33.850 62.865 ;
        RECT 33.650 62.195 33.880 62.845 ;
        RECT 34.135 62.435 34.305 63.005 ;
        RECT 34.590 62.845 34.760 65.375 ;
        RECT 35.180 65.355 35.350 65.375 ;
        RECT 35.635 65.170 35.805 66.580 ;
        RECT 36.090 66.375 36.260 66.395 ;
        RECT 36.680 66.375 36.850 66.965 ;
        RECT 36.990 66.580 37.450 66.810 ;
        RECT 36.060 65.555 36.290 66.375 ;
        RECT 36.015 65.295 36.335 65.555 ;
        RECT 36.650 65.375 36.880 66.375 ;
        RECT 36.680 65.355 36.850 65.375 ;
        RECT 35.490 64.940 35.950 65.170 ;
        RECT 35.635 64.270 35.805 64.940 ;
        RECT 35.590 63.950 35.850 64.270 ;
        RECT 36.090 64.240 36.260 65.295 ;
        RECT 37.135 65.170 37.305 66.580 ;
        RECT 37.590 66.375 37.760 66.395 ;
        RECT 38.180 66.375 38.350 66.970 ;
        RECT 39.745 66.965 40.105 66.970 ;
        RECT 42.680 66.965 43.105 66.970 ;
        RECT 45.745 66.965 46.105 66.970 ;
        RECT 38.490 66.580 38.950 66.810 ;
        RECT 39.990 66.580 40.450 66.810 ;
        RECT 41.490 66.580 41.950 66.810 ;
        RECT 37.560 65.975 37.790 66.375 ;
        RECT 37.515 65.715 37.835 65.975 ;
        RECT 37.560 65.375 37.790 65.715 ;
        RECT 38.150 65.375 38.380 66.375 ;
        RECT 36.990 64.940 37.450 65.170 ;
        RECT 37.135 64.240 37.305 64.940 ;
        RECT 36.015 63.980 36.335 64.240 ;
        RECT 37.060 63.980 37.380 64.240 ;
        RECT 35.635 63.235 35.805 63.950 ;
        RECT 35.490 63.005 35.950 63.235 ;
        RECT 35.180 62.845 35.350 62.865 ;
        RECT 33.680 61.600 33.850 62.195 ;
        RECT 34.060 62.175 34.380 62.435 ;
        RECT 34.560 62.195 34.790 62.845 ;
        RECT 35.150 62.195 35.380 62.845 ;
        RECT 34.590 62.175 34.760 62.195 ;
        RECT 34.135 62.035 34.305 62.175 ;
        RECT 33.990 61.805 34.450 62.035 ;
        RECT 35.180 61.605 35.350 62.195 ;
        RECT 35.635 62.035 35.805 63.005 ;
        RECT 36.090 62.845 36.260 63.980 ;
        RECT 37.135 63.235 37.305 63.980 ;
        RECT 36.990 63.005 37.450 63.235 ;
        RECT 36.680 62.845 36.850 62.865 ;
        RECT 36.060 62.195 36.290 62.845 ;
        RECT 36.650 62.195 36.880 62.845 ;
        RECT 36.090 62.175 36.260 62.195 ;
        RECT 35.490 61.805 35.950 62.035 ;
        RECT 35.180 61.600 35.605 61.605 ;
        RECT 36.680 61.600 36.850 62.195 ;
        RECT 37.135 62.035 37.305 63.005 ;
        RECT 37.590 62.845 37.760 65.375 ;
        RECT 38.180 65.355 38.350 65.375 ;
        RECT 38.635 65.170 38.805 66.580 ;
        RECT 39.090 66.375 39.260 66.395 ;
        RECT 39.680 66.375 39.850 66.395 ;
        RECT 39.060 65.960 39.290 66.375 ;
        RECT 39.650 65.960 39.880 66.375 ;
        RECT 40.135 65.975 40.305 66.580 ;
        RECT 41.635 66.395 41.805 66.580 ;
        RECT 40.590 66.375 40.760 66.395 ;
        RECT 41.180 66.375 41.350 66.395 ;
        RECT 39.060 65.790 39.880 65.960 ;
        RECT 39.060 65.375 39.290 65.790 ;
        RECT 39.650 65.375 39.880 65.790 ;
        RECT 40.060 65.715 40.380 65.975 ;
        RECT 40.560 65.960 40.790 66.375 ;
        RECT 41.150 65.960 41.380 66.375 ;
        RECT 41.560 66.135 41.880 66.395 ;
        RECT 42.090 66.375 42.260 66.395 ;
        RECT 42.680 66.375 42.850 66.965 ;
        RECT 42.990 66.580 43.450 66.810 ;
        RECT 44.490 66.580 44.950 66.810 ;
        RECT 45.990 66.580 46.450 66.810 ;
        RECT 40.560 65.790 41.380 65.960 ;
        RECT 39.090 65.355 39.260 65.375 ;
        RECT 39.680 65.355 39.850 65.375 ;
        RECT 40.135 65.170 40.305 65.715 ;
        RECT 40.560 65.375 40.790 65.790 ;
        RECT 41.150 65.375 41.380 65.790 ;
        RECT 40.590 65.355 40.760 65.375 ;
        RECT 41.180 65.355 41.350 65.375 ;
        RECT 41.635 65.170 41.805 66.135 ;
        RECT 42.060 65.375 42.290 66.375 ;
        RECT 42.650 65.375 42.880 66.375 ;
        RECT 38.490 64.940 38.950 65.170 ;
        RECT 39.990 64.940 40.450 65.170 ;
        RECT 41.490 64.940 41.950 65.170 ;
        RECT 38.560 64.875 38.880 64.940 ;
        RECT 38.635 63.235 38.805 64.875 ;
        RECT 39.015 63.980 39.335 64.240 ;
        RECT 38.490 63.005 38.950 63.235 ;
        RECT 38.180 62.845 38.350 62.865 ;
        RECT 37.560 62.195 37.790 62.845 ;
        RECT 38.150 62.195 38.380 62.845 ;
        RECT 37.590 62.175 37.760 62.195 ;
        RECT 36.990 61.805 37.450 62.035 ;
        RECT 38.180 61.605 38.350 62.195 ;
        RECT 38.635 62.035 38.805 63.005 ;
        RECT 39.090 62.845 39.260 63.980 ;
        RECT 40.135 63.235 40.305 64.940 ;
        RECT 40.515 63.980 40.835 64.240 ;
        RECT 39.990 63.005 40.450 63.235 ;
        RECT 39.680 62.845 39.850 62.865 ;
        RECT 39.060 62.195 39.290 62.845 ;
        RECT 39.650 62.195 39.880 62.845 ;
        RECT 39.090 62.175 39.260 62.195 ;
        RECT 38.490 61.805 38.950 62.035 ;
        RECT 38.180 61.600 38.605 61.605 ;
        RECT 39.680 61.600 39.850 62.195 ;
        RECT 40.135 62.035 40.305 63.005 ;
        RECT 40.590 62.845 40.760 63.980 ;
        RECT 41.635 63.235 41.805 64.940 ;
        RECT 42.090 64.240 42.260 65.375 ;
        RECT 42.680 65.355 42.850 65.375 ;
        RECT 43.135 65.170 43.305 66.580 ;
        RECT 43.590 66.375 43.760 66.395 ;
        RECT 44.180 66.375 44.350 66.395 ;
        RECT 43.560 65.960 43.790 66.375 ;
        RECT 44.150 65.960 44.380 66.375 ;
        RECT 43.560 65.790 44.380 65.960 ;
        RECT 43.560 65.375 43.790 65.790 ;
        RECT 44.150 65.375 44.380 65.790 ;
        RECT 44.635 65.555 44.805 66.580 ;
        RECT 46.135 66.395 46.305 66.580 ;
        RECT 45.090 66.375 45.260 66.395 ;
        RECT 45.680 66.375 45.850 66.395 ;
        RECT 45.060 65.960 45.290 66.375 ;
        RECT 45.650 65.960 45.880 66.375 ;
        RECT 46.060 66.135 46.380 66.395 ;
        RECT 46.590 66.375 46.760 66.395 ;
        RECT 45.060 65.790 45.880 65.960 ;
        RECT 43.590 65.355 43.760 65.375 ;
        RECT 44.180 65.355 44.350 65.375 ;
        RECT 44.560 65.170 44.880 65.555 ;
        RECT 45.060 65.375 45.290 65.790 ;
        RECT 45.650 65.375 45.880 65.790 ;
        RECT 45.090 65.355 45.260 65.375 ;
        RECT 45.680 65.355 45.850 65.375 ;
        RECT 46.135 65.170 46.305 66.135 ;
        RECT 46.560 65.375 46.790 66.375 ;
        RECT 42.990 64.940 43.450 65.170 ;
        RECT 44.490 64.940 44.950 65.170 ;
        RECT 45.990 64.940 46.450 65.170 ;
        RECT 43.060 64.875 43.380 64.940 ;
        RECT 42.015 63.980 42.335 64.240 ;
        RECT 41.490 63.005 41.950 63.235 ;
        RECT 41.180 62.845 41.350 62.865 ;
        RECT 40.560 62.195 40.790 62.845 ;
        RECT 41.150 62.195 41.380 62.845 ;
        RECT 40.590 62.175 40.760 62.195 ;
        RECT 39.990 61.805 40.450 62.035 ;
        RECT 41.180 61.605 41.350 62.195 ;
        RECT 41.635 62.035 41.805 63.005 ;
        RECT 42.090 62.845 42.260 63.980 ;
        RECT 43.135 63.235 43.305 64.875 ;
        RECT 43.515 63.980 43.835 64.240 ;
        RECT 42.990 63.005 43.450 63.235 ;
        RECT 42.680 62.845 42.850 62.865 ;
        RECT 42.060 62.195 42.290 62.845 ;
        RECT 42.650 62.195 42.880 62.845 ;
        RECT 42.090 62.175 42.260 62.195 ;
        RECT 41.490 61.805 41.950 62.035 ;
        RECT 41.180 61.600 41.605 61.605 ;
        RECT 42.680 61.600 42.850 62.195 ;
        RECT 43.135 62.035 43.305 63.005 ;
        RECT 43.590 62.845 43.760 63.980 ;
        RECT 44.635 63.235 44.805 64.940 ;
        RECT 45.015 63.980 45.335 64.240 ;
        RECT 44.490 63.005 44.950 63.235 ;
        RECT 44.180 62.845 44.350 62.865 ;
        RECT 43.560 62.195 43.790 62.845 ;
        RECT 44.150 62.195 44.380 62.845 ;
        RECT 43.590 62.175 43.760 62.195 ;
        RECT 42.990 61.805 43.450 62.035 ;
        RECT 44.180 61.605 44.350 62.195 ;
        RECT 44.635 62.035 44.805 63.005 ;
        RECT 45.090 62.845 45.260 63.980 ;
        RECT 46.135 63.235 46.305 64.940 ;
        RECT 46.590 64.240 46.760 65.375 ;
        RECT 46.515 63.980 46.835 64.240 ;
        RECT 45.990 63.005 46.450 63.235 ;
        RECT 45.680 62.845 45.850 62.865 ;
        RECT 45.060 62.195 45.290 62.845 ;
        RECT 45.650 62.195 45.880 62.845 ;
        RECT 45.090 62.175 45.260 62.195 ;
        RECT 44.490 61.805 44.950 62.035 ;
        RECT 44.180 61.600 44.605 61.605 ;
        RECT 45.680 61.600 45.850 62.195 ;
        RECT 46.135 62.035 46.305 63.005 ;
        RECT 46.590 62.845 46.760 63.980 ;
        RECT 46.560 62.195 46.790 62.845 ;
        RECT 46.590 62.175 46.760 62.195 ;
        RECT 45.990 61.805 46.450 62.035 ;
        RECT 33.470 61.310 46.970 61.600 ;
        RECT 35.245 61.305 35.605 61.310 ;
        RECT 38.245 61.305 38.605 61.310 ;
        RECT 41.245 61.305 41.605 61.310 ;
        RECT 44.245 61.305 44.605 61.310 ;
        RECT 33.745 60.550 34.105 60.555 ;
        RECT 36.745 60.550 37.105 60.555 ;
        RECT 39.745 60.550 40.105 60.555 ;
        RECT 42.745 60.550 43.105 60.555 ;
        RECT 45.745 60.550 46.105 60.555 ;
        RECT 33.470 60.260 46.970 60.550 ;
        RECT 33.680 60.255 34.105 60.260 ;
        RECT 33.680 59.665 33.850 60.255 ;
        RECT 33.990 59.870 34.450 60.100 ;
        RECT 33.650 58.665 33.880 59.665 ;
        RECT 33.680 58.645 33.850 58.665 ;
        RECT 34.135 58.460 34.305 59.870 ;
        RECT 34.590 59.665 34.760 59.685 ;
        RECT 35.180 59.665 35.350 60.260 ;
        RECT 36.680 60.255 37.105 60.260 ;
        RECT 35.490 59.870 35.950 60.100 ;
        RECT 34.560 58.665 34.790 59.665 ;
        RECT 35.150 58.665 35.380 59.665 ;
        RECT 33.990 58.230 34.450 58.460 ;
        RECT 34.135 56.525 34.305 58.230 ;
        RECT 33.990 56.295 34.450 56.525 ;
        RECT 33.680 56.135 33.850 56.155 ;
        RECT 33.650 55.485 33.880 56.135 ;
        RECT 33.680 54.890 33.850 55.485 ;
        RECT 34.135 55.325 34.305 56.295 ;
        RECT 34.590 56.135 34.760 58.665 ;
        RECT 35.180 58.645 35.350 58.665 ;
        RECT 35.635 58.460 35.805 59.870 ;
        RECT 36.090 59.665 36.260 59.685 ;
        RECT 36.680 59.665 36.850 60.255 ;
        RECT 36.990 59.870 37.450 60.100 ;
        RECT 36.060 58.665 36.290 59.665 ;
        RECT 36.650 58.665 36.880 59.665 ;
        RECT 35.490 58.230 35.950 58.460 ;
        RECT 36.090 58.375 36.260 58.665 ;
        RECT 36.680 58.645 36.850 58.665 ;
        RECT 37.135 58.460 37.305 59.870 ;
        RECT 37.590 59.665 37.760 59.685 ;
        RECT 38.180 59.665 38.350 60.260 ;
        RECT 39.745 60.255 40.105 60.260 ;
        RECT 42.680 60.255 43.105 60.260 ;
        RECT 45.745 60.255 46.105 60.260 ;
        RECT 38.490 59.870 38.950 60.100 ;
        RECT 39.990 59.870 40.450 60.100 ;
        RECT 41.490 59.870 41.950 60.100 ;
        RECT 37.560 58.665 37.790 59.665 ;
        RECT 38.150 58.665 38.380 59.665 ;
        RECT 36.420 58.375 36.740 58.420 ;
        RECT 35.635 57.560 35.805 58.230 ;
        RECT 36.090 58.205 36.740 58.375 ;
        RECT 36.990 58.230 37.450 58.460 ;
        RECT 35.590 57.240 35.850 57.560 ;
        RECT 36.090 57.530 36.260 58.205 ;
        RECT 36.420 58.160 36.740 58.205 ;
        RECT 37.135 57.530 37.305 58.230 ;
        RECT 36.015 57.270 36.335 57.530 ;
        RECT 37.060 57.270 37.380 57.530 ;
        RECT 35.635 56.525 35.805 57.240 ;
        RECT 35.490 56.295 35.950 56.525 ;
        RECT 35.180 56.135 35.350 56.155 ;
        RECT 34.560 55.485 34.790 56.135 ;
        RECT 35.150 55.485 35.380 56.135 ;
        RECT 34.590 55.465 34.760 55.485 ;
        RECT 33.990 55.095 34.450 55.325 ;
        RECT 34.135 54.890 34.305 55.095 ;
        RECT 35.180 54.895 35.350 55.485 ;
        RECT 35.635 55.325 35.805 56.295 ;
        RECT 36.090 56.135 36.260 57.270 ;
        RECT 37.135 56.525 37.305 57.270 ;
        RECT 36.990 56.295 37.450 56.525 ;
        RECT 36.680 56.135 36.850 56.155 ;
        RECT 36.060 55.485 36.290 56.135 ;
        RECT 36.650 55.485 36.880 56.135 ;
        RECT 36.090 55.465 36.260 55.485 ;
        RECT 35.490 55.095 35.950 55.325 ;
        RECT 35.180 54.890 35.605 54.895 ;
        RECT 36.680 54.890 36.850 55.485 ;
        RECT 37.135 55.325 37.305 56.295 ;
        RECT 37.590 56.135 37.760 58.665 ;
        RECT 38.180 58.645 38.350 58.665 ;
        RECT 38.635 58.460 38.805 59.870 ;
        RECT 39.090 59.665 39.260 59.685 ;
        RECT 39.680 59.665 39.850 59.685 ;
        RECT 39.060 59.250 39.290 59.665 ;
        RECT 39.650 59.250 39.880 59.665 ;
        RECT 40.135 59.265 40.305 59.870 ;
        RECT 41.635 59.685 41.805 59.870 ;
        RECT 40.590 59.665 40.760 59.685 ;
        RECT 41.180 59.665 41.350 59.685 ;
        RECT 39.060 59.080 39.880 59.250 ;
        RECT 39.060 58.665 39.290 59.080 ;
        RECT 39.650 58.665 39.880 59.080 ;
        RECT 40.060 59.005 40.380 59.265 ;
        RECT 40.560 59.250 40.790 59.665 ;
        RECT 41.150 59.250 41.380 59.665 ;
        RECT 41.560 59.425 41.880 59.685 ;
        RECT 42.090 59.665 42.260 59.685 ;
        RECT 42.680 59.665 42.850 60.255 ;
        RECT 42.990 59.870 43.450 60.100 ;
        RECT 44.490 59.870 44.950 60.100 ;
        RECT 45.990 59.870 46.450 60.100 ;
        RECT 40.560 59.080 41.380 59.250 ;
        RECT 39.090 58.645 39.260 58.665 ;
        RECT 39.680 58.645 39.850 58.665 ;
        RECT 40.135 58.460 40.305 59.005 ;
        RECT 40.560 58.665 40.790 59.080 ;
        RECT 41.150 58.665 41.380 59.080 ;
        RECT 40.590 58.645 40.760 58.665 ;
        RECT 41.180 58.645 41.350 58.665 ;
        RECT 41.635 58.460 41.805 59.425 ;
        RECT 42.060 58.665 42.290 59.665 ;
        RECT 42.650 58.665 42.880 59.665 ;
        RECT 38.490 58.230 38.950 58.460 ;
        RECT 39.990 58.230 40.450 58.460 ;
        RECT 41.490 58.230 41.950 58.460 ;
        RECT 38.560 58.165 38.880 58.230 ;
        RECT 38.635 56.525 38.805 58.165 ;
        RECT 39.015 57.270 39.335 57.530 ;
        RECT 38.490 56.295 38.950 56.525 ;
        RECT 38.180 56.135 38.350 56.155 ;
        RECT 37.560 55.725 37.790 56.135 ;
        RECT 37.515 55.465 37.835 55.725 ;
        RECT 38.150 55.485 38.380 56.135 ;
        RECT 36.990 55.095 37.450 55.325 ;
        RECT 38.180 54.895 38.350 55.485 ;
        RECT 38.635 55.325 38.805 56.295 ;
        RECT 39.090 56.135 39.260 57.270 ;
        RECT 40.135 56.525 40.305 58.230 ;
        RECT 40.515 57.270 40.835 57.530 ;
        RECT 39.990 56.295 40.450 56.525 ;
        RECT 39.680 56.135 39.850 56.155 ;
        RECT 39.060 55.485 39.290 56.135 ;
        RECT 39.650 55.485 39.880 56.135 ;
        RECT 39.090 55.465 39.260 55.485 ;
        RECT 38.490 55.095 38.950 55.325 ;
        RECT 38.180 54.890 38.605 54.895 ;
        RECT 39.680 54.890 39.850 55.485 ;
        RECT 40.135 55.325 40.305 56.295 ;
        RECT 40.590 56.135 40.760 57.270 ;
        RECT 41.635 56.525 41.805 58.230 ;
        RECT 42.090 57.530 42.260 58.665 ;
        RECT 42.680 58.645 42.850 58.665 ;
        RECT 43.135 58.460 43.305 59.870 ;
        RECT 43.590 59.665 43.760 59.685 ;
        RECT 44.180 59.665 44.350 59.685 ;
        RECT 43.560 59.250 43.790 59.665 ;
        RECT 44.150 59.250 44.380 59.665 ;
        RECT 43.560 59.080 44.380 59.250 ;
        RECT 43.560 58.665 43.790 59.080 ;
        RECT 44.150 58.665 44.380 59.080 ;
        RECT 44.635 58.845 44.805 59.870 ;
        RECT 46.135 59.685 46.305 59.870 ;
        RECT 45.090 59.665 45.260 59.685 ;
        RECT 45.680 59.665 45.850 59.685 ;
        RECT 45.060 59.250 45.290 59.665 ;
        RECT 45.650 59.250 45.880 59.665 ;
        RECT 46.060 59.425 46.380 59.685 ;
        RECT 46.590 59.665 46.760 59.685 ;
        RECT 45.060 59.080 45.880 59.250 ;
        RECT 43.590 58.645 43.760 58.665 ;
        RECT 44.180 58.645 44.350 58.665 ;
        RECT 44.560 58.460 44.880 58.845 ;
        RECT 45.060 58.665 45.290 59.080 ;
        RECT 45.650 58.665 45.880 59.080 ;
        RECT 45.090 58.645 45.260 58.665 ;
        RECT 45.680 58.645 45.850 58.665 ;
        RECT 46.135 58.460 46.305 59.425 ;
        RECT 46.560 58.665 46.790 59.665 ;
        RECT 42.990 58.230 43.450 58.460 ;
        RECT 44.490 58.230 44.950 58.460 ;
        RECT 45.990 58.230 46.450 58.460 ;
        RECT 43.060 58.165 43.380 58.230 ;
        RECT 42.015 57.270 42.335 57.530 ;
        RECT 41.490 56.295 41.950 56.525 ;
        RECT 41.180 56.135 41.350 56.155 ;
        RECT 40.560 55.485 40.790 56.135 ;
        RECT 41.150 55.485 41.380 56.135 ;
        RECT 40.590 55.465 40.760 55.485 ;
        RECT 39.990 55.095 40.450 55.325 ;
        RECT 41.180 54.895 41.350 55.485 ;
        RECT 41.635 55.325 41.805 56.295 ;
        RECT 42.090 56.135 42.260 57.270 ;
        RECT 43.135 56.525 43.305 58.165 ;
        RECT 43.515 57.270 43.835 57.530 ;
        RECT 42.990 56.295 43.450 56.525 ;
        RECT 42.680 56.135 42.850 56.155 ;
        RECT 42.060 55.485 42.290 56.135 ;
        RECT 42.650 55.485 42.880 56.135 ;
        RECT 42.090 55.465 42.260 55.485 ;
        RECT 41.490 55.095 41.950 55.325 ;
        RECT 41.180 54.890 41.605 54.895 ;
        RECT 42.680 54.890 42.850 55.485 ;
        RECT 43.135 55.325 43.305 56.295 ;
        RECT 43.590 56.135 43.760 57.270 ;
        RECT 44.635 56.525 44.805 58.230 ;
        RECT 45.015 57.270 45.335 57.530 ;
        RECT 44.490 56.295 44.950 56.525 ;
        RECT 44.180 56.135 44.350 56.155 ;
        RECT 43.560 55.485 43.790 56.135 ;
        RECT 44.150 55.485 44.380 56.135 ;
        RECT 43.590 55.465 43.760 55.485 ;
        RECT 42.990 55.095 43.450 55.325 ;
        RECT 44.180 54.895 44.350 55.485 ;
        RECT 44.635 55.325 44.805 56.295 ;
        RECT 45.090 56.135 45.260 57.270 ;
        RECT 46.135 56.525 46.305 58.230 ;
        RECT 46.590 57.530 46.760 58.665 ;
        RECT 46.515 57.270 46.835 57.530 ;
        RECT 45.990 56.295 46.450 56.525 ;
        RECT 45.680 56.135 45.850 56.155 ;
        RECT 45.060 55.485 45.290 56.135 ;
        RECT 45.650 55.485 45.880 56.135 ;
        RECT 45.090 55.465 45.260 55.485 ;
        RECT 44.490 55.095 44.950 55.325 ;
        RECT 44.180 54.890 44.605 54.895 ;
        RECT 45.680 54.890 45.850 55.485 ;
        RECT 46.135 55.325 46.305 56.295 ;
        RECT 46.590 56.135 46.760 57.270 ;
        RECT 46.560 55.485 46.790 56.135 ;
        RECT 46.590 55.465 46.760 55.485 ;
        RECT 45.990 55.095 46.450 55.325 ;
        RECT 33.470 54.600 46.970 54.890 ;
        RECT 35.245 54.595 35.605 54.600 ;
        RECT 38.245 54.595 38.605 54.600 ;
        RECT 41.245 54.595 41.605 54.600 ;
        RECT 44.245 54.595 44.605 54.600 ;
        RECT 33.745 53.840 34.105 53.845 ;
        RECT 36.745 53.840 37.105 53.845 ;
        RECT 39.745 53.840 40.105 53.845 ;
        RECT 42.745 53.840 43.105 53.845 ;
        RECT 45.745 53.840 46.105 53.845 ;
        RECT 33.470 53.550 46.970 53.840 ;
        RECT 33.680 53.545 34.105 53.550 ;
        RECT 33.680 52.955 33.850 53.545 ;
        RECT 33.990 53.160 34.450 53.390 ;
        RECT 33.650 51.955 33.880 52.955 ;
        RECT 33.680 51.935 33.850 51.955 ;
        RECT 34.135 51.750 34.305 53.160 ;
        RECT 34.515 52.715 34.835 52.975 ;
        RECT 35.180 52.955 35.350 53.550 ;
        RECT 36.680 53.545 37.105 53.550 ;
        RECT 35.490 53.160 35.950 53.390 ;
        RECT 34.560 51.955 34.790 52.715 ;
        RECT 35.150 51.955 35.380 52.955 ;
        RECT 33.990 51.520 34.450 51.750 ;
        RECT 34.135 49.815 34.305 51.520 ;
        RECT 33.990 49.585 34.450 49.815 ;
        RECT 33.680 49.425 33.850 49.445 ;
        RECT 33.650 48.775 33.880 49.425 ;
        RECT 34.135 49.015 34.305 49.585 ;
        RECT 34.590 49.425 34.760 51.955 ;
        RECT 35.180 51.935 35.350 51.955 ;
        RECT 35.635 51.750 35.805 53.160 ;
        RECT 36.090 52.955 36.260 52.975 ;
        RECT 36.680 52.955 36.850 53.545 ;
        RECT 36.990 53.160 37.450 53.390 ;
        RECT 36.060 52.135 36.290 52.955 ;
        RECT 36.015 51.875 36.335 52.135 ;
        RECT 36.650 51.955 36.880 52.955 ;
        RECT 36.680 51.935 36.850 51.955 ;
        RECT 35.490 51.520 35.950 51.750 ;
        RECT 35.635 50.850 35.805 51.520 ;
        RECT 35.590 50.530 35.850 50.850 ;
        RECT 36.090 50.820 36.260 51.875 ;
        RECT 37.135 51.750 37.305 53.160 ;
        RECT 37.590 52.955 37.760 52.975 ;
        RECT 38.180 52.955 38.350 53.550 ;
        RECT 39.745 53.545 40.105 53.550 ;
        RECT 42.680 53.545 43.105 53.550 ;
        RECT 45.745 53.545 46.105 53.550 ;
        RECT 38.490 53.160 38.950 53.390 ;
        RECT 39.990 53.160 40.450 53.390 ;
        RECT 41.490 53.160 41.950 53.390 ;
        RECT 37.560 52.555 37.790 52.955 ;
        RECT 37.515 52.295 37.835 52.555 ;
        RECT 37.560 51.955 37.790 52.295 ;
        RECT 38.150 51.955 38.380 52.955 ;
        RECT 36.990 51.520 37.450 51.750 ;
        RECT 37.135 50.820 37.305 51.520 ;
        RECT 36.015 50.560 36.335 50.820 ;
        RECT 37.060 50.560 37.380 50.820 ;
        RECT 35.635 49.815 35.805 50.530 ;
        RECT 35.490 49.585 35.950 49.815 ;
        RECT 35.180 49.425 35.350 49.445 ;
        RECT 33.680 48.180 33.850 48.775 ;
        RECT 34.060 48.755 34.380 49.015 ;
        RECT 34.560 48.775 34.790 49.425 ;
        RECT 35.150 48.775 35.380 49.425 ;
        RECT 34.590 48.755 34.760 48.775 ;
        RECT 34.135 48.615 34.305 48.755 ;
        RECT 33.990 48.385 34.450 48.615 ;
        RECT 35.180 48.185 35.350 48.775 ;
        RECT 35.635 48.615 35.805 49.585 ;
        RECT 36.090 49.425 36.260 50.560 ;
        RECT 37.135 49.815 37.305 50.560 ;
        RECT 36.990 49.585 37.450 49.815 ;
        RECT 36.680 49.425 36.850 49.445 ;
        RECT 36.060 48.775 36.290 49.425 ;
        RECT 36.650 48.775 36.880 49.425 ;
        RECT 36.090 48.755 36.260 48.775 ;
        RECT 35.490 48.385 35.950 48.615 ;
        RECT 35.180 48.180 35.605 48.185 ;
        RECT 36.680 48.180 36.850 48.775 ;
        RECT 37.135 48.615 37.305 49.585 ;
        RECT 37.590 49.425 37.760 51.955 ;
        RECT 38.180 51.935 38.350 51.955 ;
        RECT 38.635 51.750 38.805 53.160 ;
        RECT 39.090 52.955 39.260 52.975 ;
        RECT 39.680 52.955 39.850 52.975 ;
        RECT 39.060 52.540 39.290 52.955 ;
        RECT 39.650 52.540 39.880 52.955 ;
        RECT 40.135 52.555 40.305 53.160 ;
        RECT 41.635 52.975 41.805 53.160 ;
        RECT 40.590 52.955 40.760 52.975 ;
        RECT 41.180 52.955 41.350 52.975 ;
        RECT 39.060 52.370 39.880 52.540 ;
        RECT 39.060 51.955 39.290 52.370 ;
        RECT 39.650 51.955 39.880 52.370 ;
        RECT 40.060 52.295 40.380 52.555 ;
        RECT 40.560 52.540 40.790 52.955 ;
        RECT 41.150 52.540 41.380 52.955 ;
        RECT 41.560 52.715 41.880 52.975 ;
        RECT 42.090 52.955 42.260 52.975 ;
        RECT 42.680 52.955 42.850 53.545 ;
        RECT 42.990 53.160 43.450 53.390 ;
        RECT 44.490 53.160 44.950 53.390 ;
        RECT 45.990 53.160 46.450 53.390 ;
        RECT 40.560 52.370 41.380 52.540 ;
        RECT 39.090 51.935 39.260 51.955 ;
        RECT 39.680 51.935 39.850 51.955 ;
        RECT 40.135 51.750 40.305 52.295 ;
        RECT 40.560 51.955 40.790 52.370 ;
        RECT 41.150 51.955 41.380 52.370 ;
        RECT 40.590 51.935 40.760 51.955 ;
        RECT 41.180 51.935 41.350 51.955 ;
        RECT 41.635 51.750 41.805 52.715 ;
        RECT 42.060 51.955 42.290 52.955 ;
        RECT 42.650 51.955 42.880 52.955 ;
        RECT 38.490 51.520 38.950 51.750 ;
        RECT 39.990 51.520 40.450 51.750 ;
        RECT 41.490 51.520 41.950 51.750 ;
        RECT 38.560 51.455 38.880 51.520 ;
        RECT 38.635 49.815 38.805 51.455 ;
        RECT 39.015 50.560 39.335 50.820 ;
        RECT 38.490 49.585 38.950 49.815 ;
        RECT 38.180 49.425 38.350 49.445 ;
        RECT 37.560 48.775 37.790 49.425 ;
        RECT 38.150 48.775 38.380 49.425 ;
        RECT 37.590 48.755 37.760 48.775 ;
        RECT 36.990 48.385 37.450 48.615 ;
        RECT 38.180 48.185 38.350 48.775 ;
        RECT 38.635 48.615 38.805 49.585 ;
        RECT 39.090 49.425 39.260 50.560 ;
        RECT 40.135 49.815 40.305 51.520 ;
        RECT 40.515 50.560 40.835 50.820 ;
        RECT 39.990 49.585 40.450 49.815 ;
        RECT 39.680 49.425 39.850 49.445 ;
        RECT 39.060 48.775 39.290 49.425 ;
        RECT 39.650 48.775 39.880 49.425 ;
        RECT 39.090 48.755 39.260 48.775 ;
        RECT 38.490 48.385 38.950 48.615 ;
        RECT 38.180 48.180 38.605 48.185 ;
        RECT 39.680 48.180 39.850 48.775 ;
        RECT 40.135 48.615 40.305 49.585 ;
        RECT 40.590 49.425 40.760 50.560 ;
        RECT 41.635 49.815 41.805 51.520 ;
        RECT 42.090 50.820 42.260 51.955 ;
        RECT 42.680 51.935 42.850 51.955 ;
        RECT 43.135 51.750 43.305 53.160 ;
        RECT 43.590 52.955 43.760 52.975 ;
        RECT 44.180 52.955 44.350 52.975 ;
        RECT 43.560 52.540 43.790 52.955 ;
        RECT 44.150 52.540 44.380 52.955 ;
        RECT 43.560 52.370 44.380 52.540 ;
        RECT 43.560 51.955 43.790 52.370 ;
        RECT 44.150 51.955 44.380 52.370 ;
        RECT 44.635 52.135 44.805 53.160 ;
        RECT 46.135 52.975 46.305 53.160 ;
        RECT 45.090 52.955 45.260 52.975 ;
        RECT 45.680 52.955 45.850 52.975 ;
        RECT 45.060 52.540 45.290 52.955 ;
        RECT 45.650 52.540 45.880 52.955 ;
        RECT 46.060 52.715 46.380 52.975 ;
        RECT 46.590 52.955 46.760 52.975 ;
        RECT 45.060 52.370 45.880 52.540 ;
        RECT 43.590 51.935 43.760 51.955 ;
        RECT 44.180 51.935 44.350 51.955 ;
        RECT 44.560 51.750 44.880 52.135 ;
        RECT 45.060 51.955 45.290 52.370 ;
        RECT 45.650 51.955 45.880 52.370 ;
        RECT 45.090 51.935 45.260 51.955 ;
        RECT 45.680 51.935 45.850 51.955 ;
        RECT 46.135 51.750 46.305 52.715 ;
        RECT 46.560 51.955 46.790 52.955 ;
        RECT 42.990 51.520 43.450 51.750 ;
        RECT 44.490 51.520 44.950 51.750 ;
        RECT 45.990 51.520 46.450 51.750 ;
        RECT 43.060 51.455 43.380 51.520 ;
        RECT 42.015 50.560 42.335 50.820 ;
        RECT 41.490 49.585 41.950 49.815 ;
        RECT 41.180 49.425 41.350 49.445 ;
        RECT 40.560 48.775 40.790 49.425 ;
        RECT 41.150 48.775 41.380 49.425 ;
        RECT 40.590 48.755 40.760 48.775 ;
        RECT 39.990 48.385 40.450 48.615 ;
        RECT 41.180 48.185 41.350 48.775 ;
        RECT 41.635 48.615 41.805 49.585 ;
        RECT 42.090 49.425 42.260 50.560 ;
        RECT 43.135 49.815 43.305 51.455 ;
        RECT 43.515 50.560 43.835 50.820 ;
        RECT 42.990 49.585 43.450 49.815 ;
        RECT 42.680 49.425 42.850 49.445 ;
        RECT 42.060 48.775 42.290 49.425 ;
        RECT 42.650 48.775 42.880 49.425 ;
        RECT 42.090 48.755 42.260 48.775 ;
        RECT 41.490 48.385 41.950 48.615 ;
        RECT 41.180 48.180 41.605 48.185 ;
        RECT 42.680 48.180 42.850 48.775 ;
        RECT 43.135 48.615 43.305 49.585 ;
        RECT 43.590 49.425 43.760 50.560 ;
        RECT 44.635 49.815 44.805 51.520 ;
        RECT 45.015 50.560 45.335 50.820 ;
        RECT 44.490 49.585 44.950 49.815 ;
        RECT 44.180 49.425 44.350 49.445 ;
        RECT 43.560 48.775 43.790 49.425 ;
        RECT 44.150 48.775 44.380 49.425 ;
        RECT 43.590 48.755 43.760 48.775 ;
        RECT 42.990 48.385 43.450 48.615 ;
        RECT 44.180 48.185 44.350 48.775 ;
        RECT 44.635 48.615 44.805 49.585 ;
        RECT 45.090 49.425 45.260 50.560 ;
        RECT 46.135 49.815 46.305 51.520 ;
        RECT 46.590 50.820 46.760 51.955 ;
        RECT 59.730 51.740 60.030 51.910 ;
        RECT 61.390 51.740 61.690 52.535 ;
        RECT 63.050 51.740 63.350 53.160 ;
        RECT 46.515 50.560 46.835 50.820 ;
        RECT 45.990 49.585 46.450 49.815 ;
        RECT 45.680 49.425 45.850 49.445 ;
        RECT 45.060 48.775 45.290 49.425 ;
        RECT 45.650 48.775 45.880 49.425 ;
        RECT 45.090 48.755 45.260 48.775 ;
        RECT 44.490 48.385 44.950 48.615 ;
        RECT 44.180 48.180 44.605 48.185 ;
        RECT 45.680 48.180 45.850 48.775 ;
        RECT 46.135 48.615 46.305 49.585 ;
        RECT 46.590 49.425 46.760 50.560 ;
        RECT 48.940 49.610 49.190 51.715 ;
        RECT 46.560 48.775 46.790 49.425 ;
        RECT 46.590 48.755 46.760 48.775 ;
        RECT 45.990 48.385 46.450 48.615 ;
        RECT 33.470 47.890 46.970 48.180 ;
        RECT 49.745 48.130 50.045 51.740 ;
        RECT 50.550 49.580 51.730 51.740 ;
        RECT 52.210 49.580 53.390 51.740 ;
        RECT 53.870 49.580 55.050 51.740 ;
        RECT 55.530 49.580 56.710 51.740 ;
        RECT 57.190 49.580 58.370 51.740 ;
        RECT 58.850 49.580 60.030 51.740 ;
        RECT 60.510 49.580 61.690 51.740 ;
        RECT 62.170 50.080 63.350 51.740 ;
        RECT 62.140 49.580 63.350 50.080 ;
        RECT 63.830 49.580 65.010 51.740 ;
        RECT 65.490 49.580 66.670 51.740 ;
        RECT 67.150 49.580 68.330 51.740 ;
        RECT 68.810 49.580 69.160 51.740 ;
        RECT 69.690 49.610 69.940 51.715 ;
        RECT 51.430 48.755 51.730 49.580 ;
        RECT 53.090 49.050 53.390 49.580 ;
        RECT 53.720 48.755 54.020 48.785 ;
        RECT 55.450 48.765 69.250 49.055 ;
        RECT 51.430 48.455 54.050 48.755 ;
        RECT 53.720 48.425 54.020 48.455 ;
        RECT 55.910 48.375 56.370 48.605 ;
        RECT 55.540 48.170 55.770 48.175 ;
        RECT 53.090 48.130 53.390 48.160 ;
        RECT 35.245 47.885 35.605 47.890 ;
        RECT 38.245 47.885 38.605 47.890 ;
        RECT 41.245 47.885 41.605 47.890 ;
        RECT 44.245 47.885 44.605 47.890 ;
        RECT 49.745 47.830 53.420 48.130 ;
        RECT 53.090 47.800 53.390 47.830 ;
        RECT 51.960 47.530 52.650 47.560 ;
        RECT 54.480 47.530 55.170 47.560 ;
        RECT 33.470 46.840 55.170 47.530 ;
        RECT 33.680 46.835 34.105 46.840 ;
        RECT 33.680 46.245 33.850 46.835 ;
        RECT 33.990 46.450 34.450 46.680 ;
        RECT 33.650 45.245 33.880 46.245 ;
        RECT 33.680 45.225 33.850 45.245 ;
        RECT 34.135 45.040 34.305 46.450 ;
        RECT 34.590 46.245 34.760 46.265 ;
        RECT 35.180 46.245 35.350 46.840 ;
        RECT 36.680 46.835 37.105 46.840 ;
        RECT 35.490 46.450 35.950 46.680 ;
        RECT 34.560 45.245 34.790 46.245 ;
        RECT 35.150 45.245 35.380 46.245 ;
        RECT 33.990 44.810 34.450 45.040 ;
        RECT 33.055 44.270 33.375 44.530 ;
        RECT 34.135 43.105 34.305 44.810 ;
        RECT 33.990 42.875 34.450 43.105 ;
        RECT 33.680 42.715 33.850 42.735 ;
        RECT 33.650 42.065 33.880 42.715 ;
        RECT 33.680 41.470 33.850 42.065 ;
        RECT 34.135 41.905 34.305 42.875 ;
        RECT 34.590 42.715 34.760 45.245 ;
        RECT 35.180 45.225 35.350 45.245 ;
        RECT 35.635 45.040 35.805 46.450 ;
        RECT 36.090 46.245 36.260 46.265 ;
        RECT 36.680 46.245 36.850 46.835 ;
        RECT 36.990 46.450 37.450 46.680 ;
        RECT 36.060 45.245 36.290 46.245 ;
        RECT 36.650 45.245 36.880 46.245 ;
        RECT 35.490 44.810 35.950 45.040 ;
        RECT 36.090 44.955 36.260 45.245 ;
        RECT 36.680 45.225 36.850 45.245 ;
        RECT 37.135 45.040 37.305 46.450 ;
        RECT 37.590 46.245 37.760 46.265 ;
        RECT 38.180 46.245 38.350 46.840 ;
        RECT 39.745 46.835 40.105 46.840 ;
        RECT 42.680 46.835 43.105 46.840 ;
        RECT 45.745 46.835 46.105 46.840 ;
        RECT 38.490 46.450 38.950 46.680 ;
        RECT 39.990 46.450 40.450 46.680 ;
        RECT 41.490 46.450 41.950 46.680 ;
        RECT 37.560 45.245 37.790 46.245 ;
        RECT 38.150 45.245 38.380 46.245 ;
        RECT 36.420 44.955 36.740 45.000 ;
        RECT 35.635 44.140 35.805 44.810 ;
        RECT 36.090 44.785 36.740 44.955 ;
        RECT 36.990 44.810 37.450 45.040 ;
        RECT 35.590 43.820 35.850 44.140 ;
        RECT 36.090 44.110 36.260 44.785 ;
        RECT 36.420 44.740 36.740 44.785 ;
        RECT 37.135 44.110 37.305 44.810 ;
        RECT 36.015 43.850 36.335 44.110 ;
        RECT 37.060 43.850 37.380 44.110 ;
        RECT 35.635 43.105 35.805 43.820 ;
        RECT 35.490 42.875 35.950 43.105 ;
        RECT 35.180 42.715 35.350 42.735 ;
        RECT 34.560 42.065 34.790 42.715 ;
        RECT 35.150 42.065 35.380 42.715 ;
        RECT 34.590 42.045 34.760 42.065 ;
        RECT 33.990 41.675 34.450 41.905 ;
        RECT 34.135 41.470 34.305 41.675 ;
        RECT 35.180 41.475 35.350 42.065 ;
        RECT 35.635 41.905 35.805 42.875 ;
        RECT 36.090 42.715 36.260 43.850 ;
        RECT 37.135 43.105 37.305 43.850 ;
        RECT 36.990 42.875 37.450 43.105 ;
        RECT 36.680 42.715 36.850 42.735 ;
        RECT 36.060 42.065 36.290 42.715 ;
        RECT 36.650 42.065 36.880 42.715 ;
        RECT 36.090 42.045 36.260 42.065 ;
        RECT 35.490 41.675 35.950 41.905 ;
        RECT 35.180 41.470 35.605 41.475 ;
        RECT 36.680 41.470 36.850 42.065 ;
        RECT 37.135 41.905 37.305 42.875 ;
        RECT 37.590 42.715 37.760 45.245 ;
        RECT 38.180 45.225 38.350 45.245 ;
        RECT 38.635 45.040 38.805 46.450 ;
        RECT 39.090 46.245 39.260 46.265 ;
        RECT 39.680 46.245 39.850 46.265 ;
        RECT 39.060 45.830 39.290 46.245 ;
        RECT 39.650 45.830 39.880 46.245 ;
        RECT 40.135 45.845 40.305 46.450 ;
        RECT 41.635 46.265 41.805 46.450 ;
        RECT 40.590 46.245 40.760 46.265 ;
        RECT 41.180 46.245 41.350 46.265 ;
        RECT 39.060 45.660 39.880 45.830 ;
        RECT 39.060 45.245 39.290 45.660 ;
        RECT 39.650 45.245 39.880 45.660 ;
        RECT 40.060 45.585 40.380 45.845 ;
        RECT 40.560 45.830 40.790 46.245 ;
        RECT 41.150 45.830 41.380 46.245 ;
        RECT 41.560 46.005 41.880 46.265 ;
        RECT 42.090 46.245 42.260 46.265 ;
        RECT 42.680 46.245 42.850 46.835 ;
        RECT 51.960 46.810 52.650 46.840 ;
        RECT 54.480 46.810 55.170 46.840 ;
        RECT 55.540 47.170 55.860 48.170 ;
        RECT 42.990 46.450 43.450 46.680 ;
        RECT 44.490 46.450 44.950 46.680 ;
        RECT 45.990 46.450 46.450 46.680 ;
        RECT 40.560 45.660 41.380 45.830 ;
        RECT 39.090 45.225 39.260 45.245 ;
        RECT 39.680 45.225 39.850 45.245 ;
        RECT 40.135 45.040 40.305 45.585 ;
        RECT 40.560 45.245 40.790 45.660 ;
        RECT 41.150 45.245 41.380 45.660 ;
        RECT 40.590 45.225 40.760 45.245 ;
        RECT 41.180 45.225 41.350 45.245 ;
        RECT 41.635 45.040 41.805 46.005 ;
        RECT 42.060 45.245 42.290 46.245 ;
        RECT 42.650 45.245 42.880 46.245 ;
        RECT 38.490 44.810 38.950 45.040 ;
        RECT 39.990 44.810 40.450 45.040 ;
        RECT 41.490 44.810 41.950 45.040 ;
        RECT 38.560 44.745 38.880 44.810 ;
        RECT 38.635 43.105 38.805 44.745 ;
        RECT 39.015 43.850 39.335 44.110 ;
        RECT 38.490 42.875 38.950 43.105 ;
        RECT 38.180 42.715 38.350 42.735 ;
        RECT 37.560 42.305 37.790 42.715 ;
        RECT 37.515 42.045 37.835 42.305 ;
        RECT 38.150 42.065 38.380 42.715 ;
        RECT 36.990 41.675 37.450 41.905 ;
        RECT 38.180 41.475 38.350 42.065 ;
        RECT 38.635 41.905 38.805 42.875 ;
        RECT 39.090 42.715 39.260 43.850 ;
        RECT 40.135 43.105 40.305 44.810 ;
        RECT 40.515 43.850 40.835 44.110 ;
        RECT 39.990 42.875 40.450 43.105 ;
        RECT 39.680 42.715 39.850 42.735 ;
        RECT 39.060 42.065 39.290 42.715 ;
        RECT 39.650 42.065 39.880 42.715 ;
        RECT 39.090 42.045 39.260 42.065 ;
        RECT 38.490 41.675 38.950 41.905 ;
        RECT 38.180 41.470 38.605 41.475 ;
        RECT 39.680 41.470 39.850 42.065 ;
        RECT 40.135 41.905 40.305 42.875 ;
        RECT 40.590 42.715 40.760 43.850 ;
        RECT 41.635 43.105 41.805 44.810 ;
        RECT 42.090 44.110 42.260 45.245 ;
        RECT 42.680 45.225 42.850 45.245 ;
        RECT 43.135 45.040 43.305 46.450 ;
        RECT 43.590 46.245 43.760 46.265 ;
        RECT 44.180 46.245 44.350 46.265 ;
        RECT 43.560 45.830 43.790 46.245 ;
        RECT 44.150 45.830 44.380 46.245 ;
        RECT 43.560 45.660 44.380 45.830 ;
        RECT 43.560 45.245 43.790 45.660 ;
        RECT 44.150 45.245 44.380 45.660 ;
        RECT 44.635 45.425 44.805 46.450 ;
        RECT 46.135 46.265 46.305 46.450 ;
        RECT 55.540 46.425 55.770 47.170 ;
        RECT 56.025 46.980 56.255 48.375 ;
        RECT 56.510 48.170 56.740 48.765 ;
        RECT 57.290 48.375 57.750 48.605 ;
        RECT 56.420 47.170 56.740 48.170 ;
        RECT 56.920 48.170 57.150 48.175 ;
        RECT 56.920 47.170 57.240 48.170 ;
        RECT 55.910 46.720 56.370 46.980 ;
        RECT 45.090 46.245 45.260 46.265 ;
        RECT 45.680 46.245 45.850 46.265 ;
        RECT 45.060 45.830 45.290 46.245 ;
        RECT 45.650 45.830 45.880 46.245 ;
        RECT 46.060 46.005 46.380 46.265 ;
        RECT 46.590 46.245 46.760 46.265 ;
        RECT 45.060 45.660 45.880 45.830 ;
        RECT 43.590 45.225 43.760 45.245 ;
        RECT 44.180 45.225 44.350 45.245 ;
        RECT 44.560 45.040 44.880 45.425 ;
        RECT 45.060 45.245 45.290 45.660 ;
        RECT 45.650 45.245 45.880 45.660 ;
        RECT 45.090 45.225 45.260 45.245 ;
        RECT 45.680 45.225 45.850 45.245 ;
        RECT 46.135 45.040 46.305 46.005 ;
        RECT 46.560 45.245 46.790 46.245 ;
        RECT 55.540 46.195 56.370 46.425 ;
        RECT 55.540 45.990 55.770 45.995 ;
        RECT 42.990 44.810 43.450 45.040 ;
        RECT 44.490 44.810 44.950 45.040 ;
        RECT 45.990 44.810 46.450 45.040 ;
        RECT 43.060 44.745 43.380 44.810 ;
        RECT 42.015 43.850 42.335 44.110 ;
        RECT 41.490 42.875 41.950 43.105 ;
        RECT 41.180 42.715 41.350 42.735 ;
        RECT 40.560 42.065 40.790 42.715 ;
        RECT 41.150 42.065 41.380 42.715 ;
        RECT 40.590 42.045 40.760 42.065 ;
        RECT 39.990 41.675 40.450 41.905 ;
        RECT 41.180 41.475 41.350 42.065 ;
        RECT 41.635 41.905 41.805 42.875 ;
        RECT 42.090 42.715 42.260 43.850 ;
        RECT 43.135 43.105 43.305 44.745 ;
        RECT 43.515 43.850 43.835 44.110 ;
        RECT 42.990 42.875 43.450 43.105 ;
        RECT 42.680 42.715 42.850 42.735 ;
        RECT 42.060 42.065 42.290 42.715 ;
        RECT 42.650 42.065 42.880 42.715 ;
        RECT 42.090 42.045 42.260 42.065 ;
        RECT 41.490 41.675 41.950 41.905 ;
        RECT 41.180 41.470 41.605 41.475 ;
        RECT 42.680 41.470 42.850 42.065 ;
        RECT 43.135 41.905 43.305 42.875 ;
        RECT 43.590 42.715 43.760 43.850 ;
        RECT 44.635 43.105 44.805 44.810 ;
        RECT 45.015 43.850 45.335 44.110 ;
        RECT 44.490 42.875 44.950 43.105 ;
        RECT 44.180 42.715 44.350 42.735 ;
        RECT 43.560 42.065 43.790 42.715 ;
        RECT 44.150 42.065 44.380 42.715 ;
        RECT 43.590 42.045 43.760 42.065 ;
        RECT 42.990 41.675 43.450 41.905 ;
        RECT 44.180 41.475 44.350 42.065 ;
        RECT 44.635 41.905 44.805 42.875 ;
        RECT 45.090 42.715 45.260 43.850 ;
        RECT 46.135 43.105 46.305 44.810 ;
        RECT 46.590 44.110 46.760 45.245 ;
        RECT 55.540 44.990 55.860 45.990 ;
        RECT 46.515 43.850 46.835 44.110 ;
        RECT 45.990 42.875 46.450 43.105 ;
        RECT 45.680 42.715 45.850 42.735 ;
        RECT 45.060 42.065 45.290 42.715 ;
        RECT 45.650 42.065 45.880 42.715 ;
        RECT 45.090 42.045 45.260 42.065 ;
        RECT 44.490 41.675 44.950 41.905 ;
        RECT 44.180 41.470 44.605 41.475 ;
        RECT 45.680 41.470 45.850 42.065 ;
        RECT 46.135 41.905 46.305 42.875 ;
        RECT 46.590 42.715 46.760 43.850 ;
        RECT 46.560 42.065 46.790 42.715 ;
        RECT 55.540 42.460 55.770 44.990 ;
        RECT 56.025 44.830 56.255 46.195 ;
        RECT 56.510 46.175 56.770 46.495 ;
        RECT 56.920 46.425 57.150 47.170 ;
        RECT 57.405 46.980 57.635 48.375 ;
        RECT 57.890 48.170 58.120 48.765 ;
        RECT 58.670 48.375 59.130 48.605 ;
        RECT 57.800 47.170 58.120 48.170 ;
        RECT 58.300 48.170 58.530 48.175 ;
        RECT 58.300 47.170 58.620 48.170 ;
        RECT 57.290 46.720 57.750 46.980 ;
        RECT 56.920 46.195 57.750 46.425 ;
        RECT 56.510 45.990 56.740 46.175 ;
        RECT 56.420 44.990 56.740 45.990 ;
        RECT 55.910 44.510 56.370 44.830 ;
        RECT 55.910 42.605 56.370 42.865 ;
        RECT 46.590 42.045 46.760 42.065 ;
        RECT 45.990 41.675 46.450 41.905 ;
        RECT 55.540 41.810 55.860 42.460 ;
        RECT 56.025 41.650 56.255 42.605 ;
        RECT 56.510 42.460 56.740 44.990 ;
        RECT 56.420 41.810 56.740 42.460 ;
        RECT 56.920 45.990 57.150 45.995 ;
        RECT 56.920 44.990 57.240 45.990 ;
        RECT 56.920 42.460 57.150 44.990 ;
        RECT 57.405 44.830 57.635 46.195 ;
        RECT 57.890 46.175 58.150 46.495 ;
        RECT 58.300 46.425 58.530 47.170 ;
        RECT 58.785 46.980 59.015 48.375 ;
        RECT 59.270 48.170 59.500 48.765 ;
        RECT 60.050 48.375 60.510 48.605 ;
        RECT 59.180 47.170 59.500 48.170 ;
        RECT 59.680 48.170 59.910 48.175 ;
        RECT 59.680 47.170 60.000 48.170 ;
        RECT 58.670 46.720 59.130 46.980 ;
        RECT 58.300 46.195 59.130 46.425 ;
        RECT 57.890 45.990 58.120 46.175 ;
        RECT 57.800 44.990 58.120 45.990 ;
        RECT 57.290 44.510 57.750 44.830 ;
        RECT 57.290 42.605 57.750 42.865 ;
        RECT 56.920 41.810 57.240 42.460 ;
        RECT 57.405 41.650 57.635 42.605 ;
        RECT 57.890 42.460 58.120 44.990 ;
        RECT 57.800 41.810 58.120 42.460 ;
        RECT 58.300 45.990 58.530 45.995 ;
        RECT 58.300 44.990 58.620 45.990 ;
        RECT 58.300 42.460 58.530 44.990 ;
        RECT 58.785 44.830 59.015 46.195 ;
        RECT 59.270 46.175 59.530 46.495 ;
        RECT 59.680 46.425 59.910 47.170 ;
        RECT 60.165 46.980 60.395 48.375 ;
        RECT 60.650 48.170 60.880 48.765 ;
        RECT 61.430 48.375 61.890 48.605 ;
        RECT 60.560 47.170 60.880 48.170 ;
        RECT 61.060 48.170 61.290 48.175 ;
        RECT 61.060 47.170 61.380 48.170 ;
        RECT 60.050 46.720 60.510 46.980 ;
        RECT 59.680 46.195 60.510 46.425 ;
        RECT 59.270 45.990 59.500 46.175 ;
        RECT 59.180 44.990 59.500 45.990 ;
        RECT 58.670 44.510 59.130 44.830 ;
        RECT 58.670 42.605 59.130 42.865 ;
        RECT 58.300 41.810 58.620 42.460 ;
        RECT 58.785 41.650 59.015 42.605 ;
        RECT 59.270 42.460 59.500 44.990 ;
        RECT 59.180 41.810 59.500 42.460 ;
        RECT 59.680 45.990 59.910 45.995 ;
        RECT 59.680 44.990 60.000 45.990 ;
        RECT 59.680 42.460 59.910 44.990 ;
        RECT 60.165 44.830 60.395 46.195 ;
        RECT 60.650 46.175 60.910 46.495 ;
        RECT 61.060 46.425 61.290 47.170 ;
        RECT 61.545 46.980 61.775 48.375 ;
        RECT 62.030 48.170 62.260 48.765 ;
        RECT 62.810 48.375 63.270 48.605 ;
        RECT 61.940 47.170 62.260 48.170 ;
        RECT 62.440 48.170 62.670 48.175 ;
        RECT 62.440 47.170 62.760 48.170 ;
        RECT 61.430 46.720 61.890 46.980 ;
        RECT 61.060 46.195 61.890 46.425 ;
        RECT 60.650 45.990 60.880 46.175 ;
        RECT 60.560 44.990 60.880 45.990 ;
        RECT 60.050 44.510 60.510 44.830 ;
        RECT 60.050 42.605 60.510 42.865 ;
        RECT 59.680 41.810 60.000 42.460 ;
        RECT 60.165 41.650 60.395 42.605 ;
        RECT 60.650 42.460 60.880 44.990 ;
        RECT 60.560 41.810 60.880 42.460 ;
        RECT 61.060 45.990 61.290 45.995 ;
        RECT 61.060 44.990 61.380 45.990 ;
        RECT 61.060 42.460 61.290 44.990 ;
        RECT 61.545 44.830 61.775 46.195 ;
        RECT 62.030 46.175 62.290 46.495 ;
        RECT 62.440 46.425 62.670 47.170 ;
        RECT 62.925 46.980 63.155 48.375 ;
        RECT 63.410 48.170 63.640 48.765 ;
        RECT 64.190 48.375 64.650 48.605 ;
        RECT 63.320 47.170 63.640 48.170 ;
        RECT 63.820 48.170 64.050 48.175 ;
        RECT 63.820 47.170 64.140 48.170 ;
        RECT 62.810 46.720 63.270 46.980 ;
        RECT 62.440 46.195 63.270 46.425 ;
        RECT 62.030 45.990 62.260 46.175 ;
        RECT 61.940 44.990 62.260 45.990 ;
        RECT 61.430 44.510 61.890 44.830 ;
        RECT 61.430 42.605 61.890 42.865 ;
        RECT 61.060 41.810 61.380 42.460 ;
        RECT 61.545 41.650 61.775 42.605 ;
        RECT 62.030 42.460 62.260 44.990 ;
        RECT 61.940 41.810 62.260 42.460 ;
        RECT 62.440 45.990 62.670 45.995 ;
        RECT 62.440 44.990 62.760 45.990 ;
        RECT 62.440 42.460 62.670 44.990 ;
        RECT 62.925 44.830 63.155 46.195 ;
        RECT 63.410 46.175 63.670 46.495 ;
        RECT 63.820 46.425 64.050 47.170 ;
        RECT 64.305 46.980 64.535 48.375 ;
        RECT 64.790 48.170 65.020 48.765 ;
        RECT 65.570 48.375 66.030 48.605 ;
        RECT 64.700 47.170 65.020 48.170 ;
        RECT 65.200 48.170 65.430 48.175 ;
        RECT 65.200 47.170 65.520 48.170 ;
        RECT 64.190 46.720 64.650 46.980 ;
        RECT 63.820 46.195 64.650 46.425 ;
        RECT 63.410 45.990 63.640 46.175 ;
        RECT 63.320 44.990 63.640 45.990 ;
        RECT 62.810 44.510 63.270 44.830 ;
        RECT 62.810 42.605 63.270 42.865 ;
        RECT 62.440 41.810 62.760 42.460 ;
        RECT 62.925 41.650 63.155 42.605 ;
        RECT 63.410 42.460 63.640 44.990 ;
        RECT 63.320 41.810 63.640 42.460 ;
        RECT 63.820 45.990 64.050 45.995 ;
        RECT 63.820 44.990 64.140 45.990 ;
        RECT 63.820 42.460 64.050 44.990 ;
        RECT 64.305 44.830 64.535 46.195 ;
        RECT 64.790 46.175 65.050 46.495 ;
        RECT 65.200 46.425 65.430 47.170 ;
        RECT 65.685 46.980 65.915 48.375 ;
        RECT 66.170 48.170 66.400 48.765 ;
        RECT 66.950 48.375 67.410 48.605 ;
        RECT 66.080 47.170 66.400 48.170 ;
        RECT 66.580 48.170 66.810 48.175 ;
        RECT 66.580 47.170 66.900 48.170 ;
        RECT 65.570 46.720 66.030 46.980 ;
        RECT 65.200 46.195 66.030 46.425 ;
        RECT 64.790 45.990 65.020 46.175 ;
        RECT 64.700 44.990 65.020 45.990 ;
        RECT 64.190 44.510 64.650 44.830 ;
        RECT 64.190 42.605 64.650 42.865 ;
        RECT 63.820 41.810 64.140 42.460 ;
        RECT 64.305 41.650 64.535 42.605 ;
        RECT 64.790 42.460 65.020 44.990 ;
        RECT 64.700 41.810 65.020 42.460 ;
        RECT 65.200 45.990 65.430 45.995 ;
        RECT 65.200 44.990 65.520 45.990 ;
        RECT 65.200 42.460 65.430 44.990 ;
        RECT 65.685 44.830 65.915 46.195 ;
        RECT 66.170 46.175 66.430 46.495 ;
        RECT 66.580 46.425 66.810 47.170 ;
        RECT 67.065 46.980 67.295 48.375 ;
        RECT 67.550 48.170 67.780 48.765 ;
        RECT 68.330 48.375 68.790 48.605 ;
        RECT 67.460 47.170 67.780 48.170 ;
        RECT 67.960 48.170 68.190 48.175 ;
        RECT 67.960 47.170 68.280 48.170 ;
        RECT 66.950 46.720 67.410 46.980 ;
        RECT 66.580 46.195 67.410 46.425 ;
        RECT 66.170 45.990 66.400 46.175 ;
        RECT 66.080 44.990 66.400 45.990 ;
        RECT 65.570 44.510 66.030 44.830 ;
        RECT 65.570 42.605 66.030 42.865 ;
        RECT 65.200 41.810 65.520 42.460 ;
        RECT 65.685 41.650 65.915 42.605 ;
        RECT 66.170 42.460 66.400 44.990 ;
        RECT 66.080 41.810 66.400 42.460 ;
        RECT 66.580 45.990 66.810 45.995 ;
        RECT 66.580 44.990 66.900 45.990 ;
        RECT 66.580 42.460 66.810 44.990 ;
        RECT 67.065 44.830 67.295 46.195 ;
        RECT 67.550 46.175 67.810 46.495 ;
        RECT 67.960 46.425 68.190 47.170 ;
        RECT 68.445 46.980 68.675 48.375 ;
        RECT 68.930 48.170 69.160 48.765 ;
        RECT 68.840 47.170 69.160 48.170 ;
        RECT 68.330 46.720 68.790 46.980 ;
        RECT 67.960 46.195 68.790 46.425 ;
        RECT 67.550 45.990 67.780 46.175 ;
        RECT 67.460 44.990 67.780 45.990 ;
        RECT 66.950 44.510 67.410 44.830 ;
        RECT 66.950 42.605 67.410 42.865 ;
        RECT 66.580 41.810 66.900 42.460 ;
        RECT 67.065 41.650 67.295 42.605 ;
        RECT 67.550 42.460 67.780 44.990 ;
        RECT 67.460 41.810 67.780 42.460 ;
        RECT 67.960 45.990 68.190 45.995 ;
        RECT 67.960 44.990 68.280 45.990 ;
        RECT 67.960 42.460 68.190 44.990 ;
        RECT 68.445 44.830 68.675 46.195 ;
        RECT 68.930 46.175 69.190 46.495 ;
        RECT 68.930 45.990 69.160 46.175 ;
        RECT 68.840 44.990 69.160 45.990 ;
        RECT 68.330 44.510 68.790 44.830 ;
        RECT 68.330 42.605 68.790 42.865 ;
        RECT 67.960 41.810 68.280 42.460 ;
        RECT 68.445 41.650 68.675 42.605 ;
        RECT 68.930 42.460 69.160 44.990 ;
        RECT 68.840 41.810 69.160 42.460 ;
        RECT 50.580 41.470 51.270 41.500 ;
        RECT 54.480 41.470 55.170 41.500 ;
        RECT 33.470 40.780 55.170 41.470 ;
        RECT 55.910 41.420 56.370 41.650 ;
        RECT 57.290 41.420 57.750 41.650 ;
        RECT 58.670 41.420 59.130 41.650 ;
        RECT 60.050 41.420 60.510 41.650 ;
        RECT 61.430 41.420 61.890 41.650 ;
        RECT 62.810 41.420 63.270 41.650 ;
        RECT 64.190 41.420 64.650 41.650 ;
        RECT 65.570 41.420 66.030 41.650 ;
        RECT 66.950 41.420 67.410 41.650 ;
        RECT 68.330 41.420 68.790 41.650 ;
        RECT 56.025 41.110 56.370 41.420 ;
        RECT 57.405 41.110 57.750 41.420 ;
        RECT 58.785 41.110 59.130 41.420 ;
        RECT 60.165 41.110 60.510 41.420 ;
        RECT 61.545 41.110 61.890 41.420 ;
        RECT 62.925 41.110 63.270 41.420 ;
        RECT 64.305 41.110 64.650 41.420 ;
        RECT 65.685 41.110 66.030 41.420 ;
        RECT 67.065 41.110 67.410 41.420 ;
        RECT 68.445 41.110 68.790 41.420 ;
        RECT 55.910 40.880 56.370 41.110 ;
        RECT 57.290 40.880 57.750 41.110 ;
        RECT 58.670 40.880 59.130 41.110 ;
        RECT 60.050 40.880 60.510 41.110 ;
        RECT 61.430 40.880 61.890 41.110 ;
        RECT 62.810 40.880 63.270 41.110 ;
        RECT 64.190 40.880 64.650 41.110 ;
        RECT 65.570 40.880 66.030 41.110 ;
        RECT 66.950 40.880 67.410 41.110 ;
        RECT 68.330 40.880 68.790 41.110 ;
        RECT 50.580 40.750 51.270 40.780 ;
        RECT 54.480 40.750 55.170 40.780 ;
        RECT 33.745 40.420 34.105 40.425 ;
        RECT 36.745 40.420 37.105 40.425 ;
        RECT 39.745 40.420 40.105 40.425 ;
        RECT 42.745 40.420 43.105 40.425 ;
        RECT 45.745 40.420 46.105 40.425 ;
        RECT 33.470 40.360 46.970 40.420 ;
        RECT 33.130 40.190 46.970 40.360 ;
        RECT 32.285 37.560 32.605 37.820 ;
        RECT 16.005 37.445 16.355 37.475 ;
        RECT 16.005 37.095 28.980 37.445 ;
        RECT 16.005 37.065 16.355 37.095 ;
        RECT 33.130 35.595 33.300 40.190 ;
        RECT 33.470 40.130 46.970 40.190 ;
        RECT 33.680 40.125 34.105 40.130 ;
        RECT 33.680 39.535 33.850 40.125 ;
        RECT 33.990 39.740 34.450 39.970 ;
        RECT 33.650 38.535 33.880 39.535 ;
        RECT 33.680 38.515 33.850 38.535 ;
        RECT 34.135 38.330 34.305 39.740 ;
        RECT 34.515 39.295 34.835 39.555 ;
        RECT 35.180 39.535 35.350 40.130 ;
        RECT 36.680 40.125 37.105 40.130 ;
        RECT 35.490 39.740 35.950 39.970 ;
        RECT 34.560 38.535 34.790 39.295 ;
        RECT 35.150 38.535 35.380 39.535 ;
        RECT 33.990 38.100 34.450 38.330 ;
        RECT 34.135 36.395 34.305 38.100 ;
        RECT 33.990 36.165 34.450 36.395 ;
        RECT 33.680 36.005 33.850 36.025 ;
        RECT 33.055 35.335 33.375 35.595 ;
        RECT 33.650 35.355 33.880 36.005 ;
        RECT 34.135 35.595 34.305 36.165 ;
        RECT 34.590 36.005 34.760 38.535 ;
        RECT 35.180 38.515 35.350 38.535 ;
        RECT 35.635 38.330 35.805 39.740 ;
        RECT 36.090 39.535 36.260 39.555 ;
        RECT 36.680 39.535 36.850 40.125 ;
        RECT 36.990 39.740 37.450 39.970 ;
        RECT 36.060 38.715 36.290 39.535 ;
        RECT 36.015 38.455 36.335 38.715 ;
        RECT 36.650 38.535 36.880 39.535 ;
        RECT 36.680 38.515 36.850 38.535 ;
        RECT 35.490 38.100 35.950 38.330 ;
        RECT 35.635 37.430 35.805 38.100 ;
        RECT 35.590 37.110 35.850 37.430 ;
        RECT 36.090 37.400 36.260 38.455 ;
        RECT 37.135 38.330 37.305 39.740 ;
        RECT 37.590 39.535 37.760 39.555 ;
        RECT 38.180 39.535 38.350 40.130 ;
        RECT 39.745 40.125 40.105 40.130 ;
        RECT 42.680 40.125 43.105 40.130 ;
        RECT 45.745 40.125 46.105 40.130 ;
        RECT 38.490 39.740 38.950 39.970 ;
        RECT 39.990 39.740 40.450 39.970 ;
        RECT 41.490 39.740 41.950 39.970 ;
        RECT 37.560 39.135 37.790 39.535 ;
        RECT 37.515 38.875 37.835 39.135 ;
        RECT 37.560 38.535 37.790 38.875 ;
        RECT 38.150 38.535 38.380 39.535 ;
        RECT 36.990 38.100 37.450 38.330 ;
        RECT 37.135 37.400 37.305 38.100 ;
        RECT 36.015 37.140 36.335 37.400 ;
        RECT 37.060 37.140 37.380 37.400 ;
        RECT 35.635 36.395 35.805 37.110 ;
        RECT 35.490 36.165 35.950 36.395 ;
        RECT 35.180 36.005 35.350 36.025 ;
        RECT 33.680 34.760 33.850 35.355 ;
        RECT 34.060 35.335 34.380 35.595 ;
        RECT 34.560 35.355 34.790 36.005 ;
        RECT 35.150 35.355 35.380 36.005 ;
        RECT 34.590 35.335 34.760 35.355 ;
        RECT 34.135 35.195 34.305 35.335 ;
        RECT 33.990 34.965 34.450 35.195 ;
        RECT 35.180 34.765 35.350 35.355 ;
        RECT 35.635 35.195 35.805 36.165 ;
        RECT 36.090 36.005 36.260 37.140 ;
        RECT 37.135 36.395 37.305 37.140 ;
        RECT 36.990 36.165 37.450 36.395 ;
        RECT 36.680 36.005 36.850 36.025 ;
        RECT 36.060 35.355 36.290 36.005 ;
        RECT 36.650 35.355 36.880 36.005 ;
        RECT 36.090 35.335 36.260 35.355 ;
        RECT 35.490 34.965 35.950 35.195 ;
        RECT 35.180 34.760 35.605 34.765 ;
        RECT 36.680 34.760 36.850 35.355 ;
        RECT 37.135 35.195 37.305 36.165 ;
        RECT 37.590 36.005 37.760 38.535 ;
        RECT 38.180 38.515 38.350 38.535 ;
        RECT 38.635 38.330 38.805 39.740 ;
        RECT 39.090 39.535 39.260 39.555 ;
        RECT 39.680 39.535 39.850 39.555 ;
        RECT 39.060 39.120 39.290 39.535 ;
        RECT 39.650 39.120 39.880 39.535 ;
        RECT 40.135 39.135 40.305 39.740 ;
        RECT 41.635 39.555 41.805 39.740 ;
        RECT 40.590 39.535 40.760 39.555 ;
        RECT 41.180 39.535 41.350 39.555 ;
        RECT 39.060 38.950 39.880 39.120 ;
        RECT 39.060 38.535 39.290 38.950 ;
        RECT 39.650 38.535 39.880 38.950 ;
        RECT 40.060 38.875 40.380 39.135 ;
        RECT 40.560 39.120 40.790 39.535 ;
        RECT 41.150 39.120 41.380 39.535 ;
        RECT 41.560 39.295 41.880 39.555 ;
        RECT 42.090 39.535 42.260 39.555 ;
        RECT 42.680 39.535 42.850 40.125 ;
        RECT 55.540 40.070 55.860 40.720 ;
        RECT 42.990 39.740 43.450 39.970 ;
        RECT 44.490 39.740 44.950 39.970 ;
        RECT 45.990 39.740 46.450 39.970 ;
        RECT 56.025 39.910 56.255 40.880 ;
        RECT 56.420 40.070 56.740 40.720 ;
        RECT 56.920 40.070 57.240 40.720 ;
        RECT 40.560 38.950 41.380 39.120 ;
        RECT 39.090 38.515 39.260 38.535 ;
        RECT 39.680 38.515 39.850 38.535 ;
        RECT 40.135 38.330 40.305 38.875 ;
        RECT 40.560 38.535 40.790 38.950 ;
        RECT 41.150 38.535 41.380 38.950 ;
        RECT 40.590 38.515 40.760 38.535 ;
        RECT 41.180 38.515 41.350 38.535 ;
        RECT 41.635 38.330 41.805 39.295 ;
        RECT 42.060 38.535 42.290 39.535 ;
        RECT 42.650 38.535 42.880 39.535 ;
        RECT 38.490 38.100 38.950 38.330 ;
        RECT 39.990 38.100 40.450 38.330 ;
        RECT 41.490 38.100 41.950 38.330 ;
        RECT 38.560 38.035 38.880 38.100 ;
        RECT 38.635 36.395 38.805 38.035 ;
        RECT 39.015 37.140 39.335 37.400 ;
        RECT 38.490 36.165 38.950 36.395 ;
        RECT 38.180 36.005 38.350 36.025 ;
        RECT 37.560 35.355 37.790 36.005 ;
        RECT 38.150 35.355 38.380 36.005 ;
        RECT 37.590 35.335 37.760 35.355 ;
        RECT 36.990 34.965 37.450 35.195 ;
        RECT 38.180 34.765 38.350 35.355 ;
        RECT 38.635 35.195 38.805 36.165 ;
        RECT 39.090 36.005 39.260 37.140 ;
        RECT 40.135 36.395 40.305 38.100 ;
        RECT 40.515 37.140 40.835 37.400 ;
        RECT 39.990 36.165 40.450 36.395 ;
        RECT 39.680 36.005 39.850 36.025 ;
        RECT 39.060 35.355 39.290 36.005 ;
        RECT 39.650 35.355 39.880 36.005 ;
        RECT 39.090 35.335 39.260 35.355 ;
        RECT 38.490 34.965 38.950 35.195 ;
        RECT 38.180 34.760 38.605 34.765 ;
        RECT 39.680 34.760 39.850 35.355 ;
        RECT 40.135 35.195 40.305 36.165 ;
        RECT 40.590 36.005 40.760 37.140 ;
        RECT 41.635 36.395 41.805 38.100 ;
        RECT 42.090 37.400 42.260 38.535 ;
        RECT 42.680 38.515 42.850 38.535 ;
        RECT 43.135 38.330 43.305 39.740 ;
        RECT 43.590 39.535 43.760 39.555 ;
        RECT 44.180 39.535 44.350 39.555 ;
        RECT 43.560 39.120 43.790 39.535 ;
        RECT 44.150 39.120 44.380 39.535 ;
        RECT 43.560 38.950 44.380 39.120 ;
        RECT 43.560 38.535 43.790 38.950 ;
        RECT 44.150 38.535 44.380 38.950 ;
        RECT 44.635 38.715 44.805 39.740 ;
        RECT 46.135 39.555 46.305 39.740 ;
        RECT 55.910 39.680 56.370 39.910 ;
        RECT 45.090 39.535 45.260 39.555 ;
        RECT 45.680 39.535 45.850 39.555 ;
        RECT 45.060 39.120 45.290 39.535 ;
        RECT 45.650 39.120 45.880 39.535 ;
        RECT 46.060 39.295 46.380 39.555 ;
        RECT 46.590 39.535 46.760 39.555 ;
        RECT 45.060 38.950 45.880 39.120 ;
        RECT 43.590 38.515 43.760 38.535 ;
        RECT 44.180 38.515 44.350 38.535 ;
        RECT 44.560 38.330 44.880 38.715 ;
        RECT 45.060 38.535 45.290 38.950 ;
        RECT 45.650 38.535 45.880 38.950 ;
        RECT 45.090 38.515 45.260 38.535 ;
        RECT 45.680 38.515 45.850 38.535 ;
        RECT 46.135 38.330 46.305 39.295 ;
        RECT 46.560 38.535 46.790 39.535 ;
        RECT 56.510 39.475 56.740 40.070 ;
        RECT 57.405 39.910 57.635 40.880 ;
        RECT 57.800 40.070 58.120 40.720 ;
        RECT 58.300 40.070 58.620 40.720 ;
        RECT 57.290 39.680 57.750 39.910 ;
        RECT 57.890 39.475 58.120 40.070 ;
        RECT 58.785 39.910 59.015 40.880 ;
        RECT 59.180 40.070 59.500 40.720 ;
        RECT 59.680 40.070 60.000 40.720 ;
        RECT 58.670 39.680 59.130 39.910 ;
        RECT 59.270 39.475 59.500 40.070 ;
        RECT 60.165 39.910 60.395 40.880 ;
        RECT 60.560 40.070 60.880 40.720 ;
        RECT 61.060 40.070 61.380 40.720 ;
        RECT 60.050 39.680 60.510 39.910 ;
        RECT 60.650 39.475 60.880 40.070 ;
        RECT 61.545 39.910 61.775 40.880 ;
        RECT 61.940 40.070 62.260 40.720 ;
        RECT 62.440 40.070 62.760 40.720 ;
        RECT 61.430 39.680 61.890 39.910 ;
        RECT 62.030 39.475 62.260 40.070 ;
        RECT 62.925 39.910 63.155 40.880 ;
        RECT 63.320 40.070 63.640 40.720 ;
        RECT 63.820 40.070 64.140 40.720 ;
        RECT 62.810 39.680 63.270 39.910 ;
        RECT 63.410 39.475 63.640 40.070 ;
        RECT 64.305 39.910 64.535 40.880 ;
        RECT 64.700 40.070 65.020 40.720 ;
        RECT 65.200 40.070 65.520 40.720 ;
        RECT 64.190 39.680 64.650 39.910 ;
        RECT 64.790 39.475 65.020 40.070 ;
        RECT 65.685 39.910 65.915 40.880 ;
        RECT 66.080 40.070 66.400 40.720 ;
        RECT 66.580 40.070 66.900 40.720 ;
        RECT 65.570 39.680 66.030 39.910 ;
        RECT 66.170 39.475 66.400 40.070 ;
        RECT 67.065 39.910 67.295 40.880 ;
        RECT 67.460 40.070 67.780 40.720 ;
        RECT 67.960 40.070 68.280 40.720 ;
        RECT 66.950 39.680 67.410 39.910 ;
        RECT 67.550 39.475 67.780 40.070 ;
        RECT 68.445 39.910 68.675 40.880 ;
        RECT 68.840 40.070 69.160 40.720 ;
        RECT 68.330 39.680 68.790 39.910 ;
        RECT 68.930 39.475 69.160 40.070 ;
        RECT 55.450 39.185 69.250 39.475 ;
        RECT 102.225 38.950 102.575 41.110 ;
        RECT 103.055 38.950 104.235 41.110 ;
        RECT 104.715 38.950 105.895 41.110 ;
        RECT 106.375 38.950 107.555 41.110 ;
        RECT 108.035 38.950 109.215 41.110 ;
        RECT 109.695 38.950 110.875 41.110 ;
        RECT 111.355 38.950 112.535 41.110 ;
        RECT 113.015 38.950 114.195 41.110 ;
        RECT 114.675 38.950 115.855 41.110 ;
        RECT 116.335 38.950 117.515 41.110 ;
        RECT 117.995 38.950 119.175 41.110 ;
        RECT 119.655 38.950 120.835 41.110 ;
        RECT 121.315 38.950 121.665 41.110 ;
        RECT 42.990 38.100 43.450 38.330 ;
        RECT 44.490 38.100 44.950 38.330 ;
        RECT 45.990 38.100 46.450 38.330 ;
        RECT 43.060 38.035 43.380 38.100 ;
        RECT 42.015 37.140 42.335 37.400 ;
        RECT 41.490 36.165 41.950 36.395 ;
        RECT 41.180 36.005 41.350 36.025 ;
        RECT 40.560 35.355 40.790 36.005 ;
        RECT 41.150 35.355 41.380 36.005 ;
        RECT 40.590 35.335 40.760 35.355 ;
        RECT 39.990 34.965 40.450 35.195 ;
        RECT 41.180 34.765 41.350 35.355 ;
        RECT 41.635 35.195 41.805 36.165 ;
        RECT 42.090 36.005 42.260 37.140 ;
        RECT 43.135 36.395 43.305 38.035 ;
        RECT 43.515 37.140 43.835 37.400 ;
        RECT 42.990 36.165 43.450 36.395 ;
        RECT 42.680 36.005 42.850 36.025 ;
        RECT 42.060 35.355 42.290 36.005 ;
        RECT 42.650 35.355 42.880 36.005 ;
        RECT 42.090 35.335 42.260 35.355 ;
        RECT 41.490 34.965 41.950 35.195 ;
        RECT 41.180 34.760 41.605 34.765 ;
        RECT 42.680 34.760 42.850 35.355 ;
        RECT 43.135 35.195 43.305 36.165 ;
        RECT 43.590 36.005 43.760 37.140 ;
        RECT 44.635 36.395 44.805 38.100 ;
        RECT 45.015 37.140 45.335 37.400 ;
        RECT 44.490 36.165 44.950 36.395 ;
        RECT 44.180 36.005 44.350 36.025 ;
        RECT 43.560 35.355 43.790 36.005 ;
        RECT 44.150 35.355 44.380 36.005 ;
        RECT 43.590 35.335 43.760 35.355 ;
        RECT 42.990 34.965 43.450 35.195 ;
        RECT 44.180 34.765 44.350 35.355 ;
        RECT 44.635 35.195 44.805 36.165 ;
        RECT 45.090 36.005 45.260 37.140 ;
        RECT 46.135 36.395 46.305 38.100 ;
        RECT 46.590 37.400 46.760 38.535 ;
        RECT 57.230 38.420 65.080 38.610 ;
        RECT 56.000 37.835 56.960 38.155 ;
        RECT 57.230 38.035 57.560 38.420 ;
        RECT 57.880 37.835 58.840 38.155 ;
        RECT 59.110 38.035 59.440 38.420 ;
        RECT 59.760 37.875 60.720 38.205 ;
        RECT 60.990 38.035 61.320 38.420 ;
        RECT 61.640 38.105 62.600 38.205 ;
        RECT 61.640 37.895 62.730 38.105 ;
        RECT 62.870 38.035 63.200 38.420 ;
        RECT 61.640 37.875 62.850 37.895 ;
        RECT 63.520 37.880 64.480 38.110 ;
        RECT 64.750 38.035 65.080 38.420 ;
        RECT 65.400 38.105 66.360 38.110 ;
        RECT 65.400 37.880 66.640 38.105 ;
        RECT 46.515 37.140 46.835 37.400 ;
        RECT 45.990 36.165 46.450 36.395 ;
        RECT 45.680 36.005 45.850 36.025 ;
        RECT 45.060 35.355 45.290 36.005 ;
        RECT 45.650 35.355 45.880 36.005 ;
        RECT 45.090 35.335 45.260 35.355 ;
        RECT 44.490 34.965 44.950 35.195 ;
        RECT 44.180 34.760 44.605 34.765 ;
        RECT 45.680 34.760 45.850 35.355 ;
        RECT 46.135 35.195 46.305 36.165 ;
        RECT 46.590 36.005 46.760 37.140 ;
        RECT 46.560 35.355 46.790 36.005 ;
        RECT 46.590 35.335 46.760 35.355 ;
        RECT 45.990 34.965 46.450 35.195 ;
        RECT 33.470 34.470 46.970 34.760 ;
        RECT 35.245 34.465 35.605 34.470 ;
        RECT 38.245 34.465 38.605 34.470 ;
        RECT 41.245 34.465 41.605 34.470 ;
        RECT 44.245 34.465 44.605 34.470 ;
        RECT 55.720 33.915 55.950 37.675 ;
        RECT 55.635 33.675 55.950 33.915 ;
        RECT 55.635 32.495 55.825 33.675 ;
        RECT 56.385 33.470 56.575 37.835 ;
        RECT 57.010 37.625 57.240 37.675 ;
        RECT 57.600 37.625 57.830 37.675 ;
        RECT 57.010 37.435 57.830 37.625 ;
        RECT 57.010 33.915 57.240 37.435 ;
        RECT 57.010 33.910 57.355 33.915 ;
        RECT 57.600 33.910 57.830 37.435 ;
        RECT 57.010 33.675 57.830 33.910 ;
        RECT 56.000 33.240 56.960 33.470 ;
        RECT 56.060 32.930 56.900 33.240 ;
        RECT 57.165 33.175 57.705 33.675 ;
        RECT 58.265 33.470 58.455 37.835 ;
        RECT 58.890 33.920 59.120 37.675 ;
        RECT 58.890 33.675 59.205 33.920 ;
        RECT 59.480 33.915 59.710 37.675 ;
        RECT 57.880 33.240 58.840 33.470 ;
        RECT 57.155 32.985 57.705 33.175 ;
        RECT 56.000 32.700 56.960 32.930 ;
        RECT 55.635 32.250 55.950 32.495 ;
        RECT 55.720 29.095 55.950 32.250 ;
        RECT 55.580 28.495 56.180 29.095 ;
        RECT 55.580 27.345 55.775 28.495 ;
        RECT 56.385 28.290 56.575 32.700 ;
        RECT 57.165 32.495 57.705 32.985 ;
        RECT 57.890 32.930 58.830 33.240 ;
        RECT 57.880 32.700 58.840 32.930 ;
        RECT 57.010 32.255 57.830 32.495 ;
        RECT 57.010 32.250 57.355 32.255 ;
        RECT 57.010 28.735 57.240 32.250 ;
        RECT 57.600 28.735 57.830 32.255 ;
        RECT 57.010 28.545 57.830 28.735 ;
        RECT 57.010 28.495 57.240 28.545 ;
        RECT 57.600 28.495 57.830 28.545 ;
        RECT 58.265 28.290 58.455 32.700 ;
        RECT 59.015 32.495 59.205 33.675 ;
        RECT 58.890 32.260 59.205 32.495 ;
        RECT 59.375 33.675 59.710 33.915 ;
        RECT 59.375 32.495 59.565 33.675 ;
        RECT 60.145 33.475 60.335 37.875 ;
        RECT 62.025 37.675 62.850 37.875 ;
        RECT 60.770 37.135 61.590 37.675 ;
        RECT 60.770 33.915 61.000 37.135 ;
        RECT 61.360 33.915 61.590 37.135 ;
        RECT 60.770 33.675 61.590 33.915 ;
        RECT 62.025 37.445 62.880 37.675 ;
        RECT 62.025 33.925 62.215 37.445 ;
        RECT 62.650 33.925 62.880 37.445 ;
        RECT 63.150 37.085 63.750 37.685 ;
        RECT 62.025 33.920 62.960 33.925 ;
        RECT 59.760 32.695 60.720 33.475 ;
        RECT 59.375 32.260 59.710 32.495 ;
        RECT 58.890 28.740 59.120 32.260 ;
        RECT 59.480 29.105 59.710 32.260 ;
        RECT 58.890 28.495 59.205 28.740 ;
        RECT 56.000 28.060 56.960 28.290 ;
        RECT 57.880 28.060 58.840 28.290 ;
        RECT 59.015 27.735 59.205 28.495 ;
        RECT 56.000 27.715 56.960 27.735 ;
        RECT 57.880 27.715 59.205 27.735 ;
        RECT 56.000 27.525 59.205 27.715 ;
        RECT 56.000 27.505 56.960 27.525 ;
        RECT 57.880 27.505 59.205 27.525 ;
        RECT 55.580 26.735 56.180 27.345 ;
        RECT 55.720 25.585 55.950 26.735 ;
        RECT 55.635 25.345 55.950 25.585 ;
        RECT 55.635 24.255 55.825 25.345 ;
        RECT 56.385 25.185 56.575 27.505 ;
        RECT 57.010 27.295 57.240 27.345 ;
        RECT 57.600 27.295 57.830 27.345 ;
        RECT 57.010 27.105 57.830 27.295 ;
        RECT 57.010 25.585 57.240 27.105 ;
        RECT 57.600 25.585 57.830 27.105 ;
        RECT 58.260 27.100 59.205 27.505 ;
        RECT 59.380 28.505 59.990 29.105 ;
        RECT 59.380 28.495 59.710 28.505 ;
        RECT 59.380 27.345 59.570 28.495 ;
        RECT 60.145 28.290 60.335 32.695 ;
        RECT 60.905 32.495 61.465 33.675 ;
        RECT 62.025 33.475 62.965 33.920 ;
        RECT 63.240 33.915 63.470 37.085 ;
        RECT 61.640 32.695 62.965 33.475 ;
        RECT 60.770 32.245 61.590 32.495 ;
        RECT 62.020 32.265 62.965 32.695 ;
        RECT 60.770 28.735 61.000 32.245 ;
        RECT 61.360 28.735 61.590 32.245 ;
        RECT 60.770 28.545 61.590 28.735 ;
        RECT 62.025 32.260 62.965 32.265 ;
        RECT 63.145 33.675 63.470 33.915 ;
        RECT 63.145 32.495 63.335 33.675 ;
        RECT 63.905 33.475 64.095 37.880 ;
        RECT 64.530 33.915 64.760 37.675 ;
        RECT 65.040 37.085 65.640 37.685 ;
        RECT 65.780 37.445 66.640 37.880 ;
        RECT 65.120 33.930 65.350 37.085 ;
        RECT 64.530 33.675 64.845 33.915 ;
        RECT 63.500 32.695 64.500 33.475 ;
        RECT 63.145 32.260 63.470 32.495 ;
        RECT 62.025 32.255 62.960 32.260 ;
        RECT 62.025 28.725 62.215 32.255 ;
        RECT 62.650 28.735 62.880 32.255 ;
        RECT 62.650 28.725 62.975 28.735 ;
        RECT 60.770 28.495 61.000 28.545 ;
        RECT 61.360 28.495 61.590 28.545 ;
        RECT 62.020 28.290 62.975 28.725 ;
        RECT 63.240 28.495 63.470 32.260 ;
        RECT 63.905 28.290 64.095 32.695 ;
        RECT 64.655 32.495 64.845 33.675 ;
        RECT 64.530 32.290 64.845 32.495 ;
        RECT 65.025 33.675 65.350 33.930 ;
        RECT 65.785 33.915 65.975 37.445 ;
        RECT 66.410 33.920 66.640 37.445 ;
        RECT 67.140 36.515 68.330 38.675 ;
        RECT 68.800 36.515 69.990 38.675 ;
        RECT 102.225 36.515 103.415 38.675 ;
        RECT 103.885 36.515 105.075 38.675 ;
        RECT 107.135 38.420 114.985 38.610 ;
        RECT 105.855 38.105 106.815 38.110 ;
        RECT 105.575 37.880 106.815 38.105 ;
        RECT 107.135 38.035 107.465 38.420 ;
        RECT 107.735 37.880 108.695 38.110 ;
        RECT 109.015 38.035 109.345 38.420 ;
        RECT 109.615 38.105 110.575 38.205 ;
        RECT 109.485 37.895 110.575 38.105 ;
        RECT 110.895 38.035 111.225 38.420 ;
        RECT 105.575 37.445 106.435 37.880 ;
        RECT 105.575 33.920 105.805 37.445 ;
        RECT 66.410 33.915 66.725 33.920 ;
        RECT 65.025 32.495 65.215 33.675 ;
        RECT 65.785 33.475 66.725 33.915 ;
        RECT 65.380 32.695 66.725 33.475 ;
        RECT 64.530 29.035 64.760 32.290 ;
        RECT 65.025 32.270 65.350 32.495 ;
        RECT 64.340 28.435 64.950 29.035 ;
        RECT 65.120 28.495 65.350 32.270 ;
        RECT 65.785 32.255 66.725 32.695 ;
        RECT 65.785 28.725 65.975 32.255 ;
        RECT 66.410 32.250 66.725 32.255 ;
        RECT 105.490 33.915 105.805 33.920 ;
        RECT 106.240 33.915 106.430 37.445 ;
        RECT 106.575 37.085 107.175 37.685 ;
        RECT 105.490 33.475 106.430 33.915 ;
        RECT 106.865 33.930 107.095 37.085 ;
        RECT 106.865 33.675 107.190 33.930 ;
        RECT 107.455 33.915 107.685 37.675 ;
        RECT 105.490 32.695 106.835 33.475 ;
        RECT 105.490 32.255 106.430 32.695 ;
        RECT 107.000 32.495 107.190 33.675 ;
        RECT 105.490 32.250 105.805 32.255 ;
        RECT 66.410 29.035 66.640 32.250 ;
        RECT 86.170 31.835 87.550 32.125 ;
        RECT 86.630 31.445 87.090 31.675 ;
        RECT 86.260 31.240 86.490 31.245 ;
        RECT 66.220 28.725 66.830 29.035 ;
        RECT 65.780 28.435 66.830 28.725 ;
        RECT 65.780 28.290 66.610 28.435 ;
        RECT 59.760 28.285 60.720 28.290 ;
        RECT 61.640 28.285 62.975 28.290 ;
        RECT 59.760 28.055 62.975 28.285 ;
        RECT 63.520 28.060 64.480 28.290 ;
        RECT 65.400 28.095 66.610 28.290 ;
        RECT 65.400 28.060 66.360 28.095 ;
        RECT 59.760 27.505 60.720 27.735 ;
        RECT 61.640 27.505 62.600 27.735 ;
        RECT 59.380 27.335 59.710 27.345 ;
        RECT 58.260 27.095 59.200 27.100 ;
        RECT 57.010 25.345 57.830 25.585 ;
        RECT 58.265 25.585 58.455 27.095 ;
        RECT 58.890 25.585 59.120 27.095 ;
        RECT 59.380 26.735 59.990 27.335 ;
        RECT 59.480 25.585 59.710 26.735 ;
        RECT 56.000 24.415 56.960 25.185 ;
        RECT 55.635 24.020 55.950 24.255 ;
        RECT 55.720 22.255 55.950 24.020 ;
        RECT 56.385 22.135 56.575 24.415 ;
        RECT 57.130 24.255 57.695 25.345 ;
        RECT 58.265 25.195 59.215 25.585 ;
        RECT 57.880 24.415 59.215 25.195 ;
        RECT 57.010 24.005 57.830 24.255 ;
        RECT 57.010 22.885 57.240 24.005 ;
        RECT 57.600 22.885 57.830 24.005 ;
        RECT 57.010 22.285 57.830 22.885 ;
        RECT 58.265 24.015 59.215 24.415 ;
        RECT 58.265 22.485 58.455 24.015 ;
        RECT 58.890 24.010 59.215 24.015 ;
        RECT 59.395 25.345 59.710 25.585 ;
        RECT 59.395 24.255 59.585 25.345 ;
        RECT 60.145 25.185 60.335 27.505 ;
        RECT 60.770 27.295 61.000 27.345 ;
        RECT 61.360 27.295 61.590 27.345 ;
        RECT 60.770 27.105 61.590 27.295 ;
        RECT 60.770 25.585 61.000 27.105 ;
        RECT 61.360 25.585 61.590 27.105 ;
        RECT 60.770 25.345 61.590 25.585 ;
        RECT 59.760 24.415 60.720 25.185 ;
        RECT 58.890 22.485 59.120 24.010 ;
        RECT 59.395 24.000 59.710 24.255 ;
        RECT 57.010 22.255 57.240 22.285 ;
        RECT 57.600 22.255 57.830 22.285 ;
        RECT 58.260 22.255 59.120 22.485 ;
        RECT 59.480 22.255 59.710 24.000 ;
        RECT 58.260 22.135 59.100 22.255 ;
        RECT 56.030 22.095 56.930 22.135 ;
        RECT 57.910 22.095 59.100 22.135 ;
        RECT 60.145 22.095 60.335 24.415 ;
        RECT 60.905 24.255 61.465 25.345 ;
        RECT 62.025 25.185 62.215 27.505 ;
        RECT 62.785 27.345 62.975 28.055 ;
        RECT 67.200 27.735 67.450 30.400 ;
        RECT 67.970 28.265 69.160 30.425 ;
        RECT 69.640 28.235 69.990 30.455 ;
        RECT 86.260 30.240 86.580 31.240 ;
        RECT 86.260 29.495 86.490 30.240 ;
        RECT 86.745 30.050 86.975 31.445 ;
        RECT 87.230 31.240 87.460 31.835 ;
        RECT 87.140 30.240 87.460 31.240 ;
        RECT 86.630 29.790 87.090 30.050 ;
        RECT 86.260 29.265 87.090 29.495 ;
        RECT 86.260 29.060 86.490 29.065 ;
        RECT 86.260 28.060 86.580 29.060 ;
        RECT 63.500 27.505 68.520 27.735 ;
        RECT 62.650 27.100 62.975 27.345 ;
        RECT 62.650 25.590 62.880 27.100 ;
        RECT 62.650 25.345 62.965 25.590 ;
        RECT 63.240 25.585 63.470 27.345 ;
        RECT 61.640 24.415 62.600 25.185 ;
        RECT 60.770 24.015 61.590 24.255 ;
        RECT 60.770 22.495 61.000 24.015 ;
        RECT 61.360 22.495 61.590 24.015 ;
        RECT 60.770 22.305 61.590 22.495 ;
        RECT 60.770 22.255 61.000 22.305 ;
        RECT 61.360 22.255 61.590 22.305 ;
        RECT 62.025 22.095 62.215 24.415 ;
        RECT 62.775 24.255 62.965 25.345 ;
        RECT 62.650 24.015 62.965 24.255 ;
        RECT 63.155 25.345 63.470 25.585 ;
        RECT 63.155 24.255 63.345 25.345 ;
        RECT 63.905 25.185 64.095 27.505 ;
        RECT 64.530 27.335 64.760 27.345 ;
        RECT 64.350 26.735 64.950 27.335 ;
        RECT 64.530 25.590 64.760 26.735 ;
        RECT 64.530 25.345 64.845 25.590 ;
        RECT 65.120 25.585 65.350 27.345 ;
        RECT 63.500 24.415 64.500 25.185 ;
        RECT 62.650 22.255 62.880 24.015 ;
        RECT 63.155 24.010 63.470 24.255 ;
        RECT 63.240 22.855 63.470 24.010 ;
        RECT 63.160 22.255 63.760 22.855 ;
        RECT 63.905 22.095 64.095 24.415 ;
        RECT 64.655 24.255 64.845 25.345 ;
        RECT 64.530 24.010 64.845 24.255 ;
        RECT 65.025 25.345 65.350 25.585 ;
        RECT 65.025 24.255 65.215 25.345 ;
        RECT 65.785 25.185 65.975 27.505 ;
        RECT 66.410 27.335 66.640 27.345 ;
        RECT 66.230 26.735 66.830 27.335 ;
        RECT 66.410 25.585 66.640 26.735 ;
        RECT 67.000 25.590 67.230 27.345 ;
        RECT 66.410 25.345 66.725 25.585 ;
        RECT 65.380 24.415 66.380 25.185 ;
        RECT 64.530 22.255 64.760 24.010 ;
        RECT 65.025 24.000 65.350 24.255 ;
        RECT 65.120 22.855 65.350 24.000 ;
        RECT 65.040 22.255 65.640 22.855 ;
        RECT 65.785 22.095 65.975 24.415 ;
        RECT 66.535 24.255 66.725 25.345 ;
        RECT 66.410 24.000 66.725 24.255 ;
        RECT 66.905 25.345 67.230 25.590 ;
        RECT 67.660 27.115 68.520 27.505 ;
        RECT 67.660 25.595 67.855 27.115 ;
        RECT 68.290 25.595 68.520 27.115 ;
        RECT 69.720 26.865 69.990 26.955 ;
        RECT 68.765 26.675 69.990 26.865 ;
        RECT 67.660 25.590 68.610 25.595 ;
        RECT 66.905 24.255 67.095 25.345 ;
        RECT 67.660 25.185 68.615 25.590 ;
        RECT 67.260 24.415 68.615 25.185 ;
        RECT 66.905 24.000 67.230 24.255 ;
        RECT 66.410 22.255 66.640 24.000 ;
        RECT 67.000 22.855 67.230 24.000 ;
        RECT 67.660 24.025 68.615 24.415 ;
        RECT 66.920 22.255 67.520 22.855 ;
        RECT 67.660 22.495 67.855 24.025 ;
        RECT 68.290 24.015 68.615 24.025 ;
        RECT 68.765 25.580 68.955 26.675 ;
        RECT 69.720 26.575 69.990 26.675 ;
        RECT 69.760 26.540 69.950 26.575 ;
        RECT 69.720 25.580 69.990 25.670 ;
        RECT 68.765 25.390 69.990 25.580 ;
        RECT 68.765 24.295 68.955 25.390 ;
        RECT 69.720 25.290 69.990 25.390 ;
        RECT 86.260 25.530 86.490 28.060 ;
        RECT 86.745 27.900 86.975 29.265 ;
        RECT 87.230 29.245 87.490 29.565 ;
        RECT 87.230 29.060 87.460 29.245 ;
        RECT 87.140 28.060 87.460 29.060 ;
        RECT 102.225 28.235 102.575 30.455 ;
        RECT 103.055 28.265 104.245 30.425 ;
        RECT 86.630 27.580 87.090 27.900 ;
        RECT 86.630 25.675 87.090 25.935 ;
        RECT 69.760 25.260 69.950 25.290 ;
        RECT 86.260 24.880 86.580 25.530 ;
        RECT 86.745 24.720 86.975 25.675 ;
        RECT 87.230 25.530 87.460 28.060 ;
        RECT 104.765 27.735 105.015 30.400 ;
        RECT 105.575 29.035 105.805 32.250 ;
        RECT 105.385 28.725 105.995 29.035 ;
        RECT 106.240 28.725 106.430 32.255 ;
        RECT 106.865 32.270 107.190 32.495 ;
        RECT 107.370 33.675 107.685 33.915 ;
        RECT 107.370 32.495 107.560 33.675 ;
        RECT 108.120 33.475 108.310 37.880 ;
        RECT 109.365 37.875 110.575 37.895 ;
        RECT 111.495 37.875 112.455 38.205 ;
        RECT 112.775 38.035 113.105 38.420 ;
        RECT 108.465 37.085 109.065 37.685 ;
        RECT 109.365 37.675 110.190 37.875 ;
        RECT 109.335 37.445 110.190 37.675 ;
        RECT 108.745 33.915 108.975 37.085 ;
        RECT 109.335 33.925 109.565 37.445 ;
        RECT 110.000 33.925 110.190 37.445 ;
        RECT 109.255 33.920 110.190 33.925 ;
        RECT 108.745 33.675 109.070 33.915 ;
        RECT 107.715 32.695 108.715 33.475 ;
        RECT 107.370 32.290 107.685 32.495 ;
        RECT 105.385 28.435 106.435 28.725 ;
        RECT 106.865 28.495 107.095 32.270 ;
        RECT 107.455 29.035 107.685 32.290 ;
        RECT 107.265 28.435 107.875 29.035 ;
        RECT 105.605 28.290 106.435 28.435 ;
        RECT 108.120 28.290 108.310 32.695 ;
        RECT 108.880 32.495 109.070 33.675 ;
        RECT 108.745 32.260 109.070 32.495 ;
        RECT 109.250 33.475 110.190 33.920 ;
        RECT 110.625 37.135 111.445 37.675 ;
        RECT 110.625 33.915 110.855 37.135 ;
        RECT 111.215 33.915 111.445 37.135 ;
        RECT 110.625 33.675 111.445 33.915 ;
        RECT 109.250 32.695 110.575 33.475 ;
        RECT 109.250 32.265 110.195 32.695 ;
        RECT 110.750 32.495 111.310 33.675 ;
        RECT 111.880 33.475 112.070 37.875 ;
        RECT 113.375 37.835 114.335 38.155 ;
        RECT 114.655 38.035 114.985 38.420 ;
        RECT 115.255 37.835 116.215 38.155 ;
        RECT 112.505 33.915 112.735 37.675 ;
        RECT 113.095 33.920 113.325 37.675 ;
        RECT 112.505 33.675 112.840 33.915 ;
        RECT 111.495 32.695 112.455 33.475 ;
        RECT 109.250 32.260 110.190 32.265 ;
        RECT 108.745 28.495 108.975 32.260 ;
        RECT 109.255 32.255 110.190 32.260 ;
        RECT 109.335 28.735 109.565 32.255 ;
        RECT 109.240 28.725 109.565 28.735 ;
        RECT 110.000 28.725 110.190 32.255 ;
        RECT 110.625 32.245 111.445 32.495 ;
        RECT 110.625 28.735 110.855 32.245 ;
        RECT 111.215 28.735 111.445 32.245 ;
        RECT 109.240 28.290 110.195 28.725 ;
        RECT 110.625 28.545 111.445 28.735 ;
        RECT 110.625 28.495 110.855 28.545 ;
        RECT 111.215 28.495 111.445 28.545 ;
        RECT 111.880 28.290 112.070 32.695 ;
        RECT 112.650 32.495 112.840 33.675 ;
        RECT 112.505 32.260 112.840 32.495 ;
        RECT 113.010 33.675 113.325 33.920 ;
        RECT 113.010 32.495 113.200 33.675 ;
        RECT 113.760 33.470 113.950 37.835 ;
        RECT 114.385 37.625 114.615 37.675 ;
        RECT 114.975 37.625 115.205 37.675 ;
        RECT 114.385 37.435 115.205 37.625 ;
        RECT 114.385 33.910 114.615 37.435 ;
        RECT 114.975 33.915 115.205 37.435 ;
        RECT 114.860 33.910 115.205 33.915 ;
        RECT 114.385 33.675 115.205 33.910 ;
        RECT 113.375 33.240 114.335 33.470 ;
        RECT 113.385 32.930 114.325 33.240 ;
        RECT 114.510 33.175 115.050 33.675 ;
        RECT 115.640 33.470 115.830 37.835 ;
        RECT 116.265 33.915 116.495 37.675 ;
        RECT 116.265 33.675 116.580 33.915 ;
        RECT 115.255 33.240 116.215 33.470 ;
        RECT 114.510 32.985 115.060 33.175 ;
        RECT 113.375 32.700 114.335 32.930 ;
        RECT 113.010 32.260 113.325 32.495 ;
        RECT 112.505 29.105 112.735 32.260 ;
        RECT 112.225 28.505 112.835 29.105 ;
        RECT 113.095 28.740 113.325 32.260 ;
        RECT 112.505 28.495 112.835 28.505 ;
        RECT 105.605 28.095 106.815 28.290 ;
        RECT 105.855 28.060 106.815 28.095 ;
        RECT 107.735 28.060 108.695 28.290 ;
        RECT 109.240 28.285 110.575 28.290 ;
        RECT 111.495 28.285 112.455 28.290 ;
        RECT 109.240 28.055 112.455 28.285 ;
        RECT 103.695 27.505 108.715 27.735 ;
        RECT 103.695 27.115 104.555 27.505 ;
        RECT 102.225 26.865 102.495 26.955 ;
        RECT 102.225 26.675 103.450 26.865 ;
        RECT 102.225 26.575 102.495 26.675 ;
        RECT 102.265 26.540 102.455 26.575 ;
        RECT 87.140 24.880 87.460 25.530 ;
        RECT 102.225 25.580 102.495 25.670 ;
        RECT 103.260 25.580 103.450 26.675 ;
        RECT 103.695 25.595 103.925 27.115 ;
        RECT 104.360 25.595 104.555 27.115 ;
        RECT 103.605 25.590 104.555 25.595 ;
        RECT 102.225 25.390 103.450 25.580 ;
        RECT 102.225 25.290 102.495 25.390 ;
        RECT 102.265 25.260 102.455 25.290 ;
        RECT 86.630 24.490 87.090 24.720 ;
        RECT 69.720 24.295 69.990 24.385 ;
        RECT 68.765 24.105 69.990 24.295 ;
        RECT 86.745 24.180 87.090 24.490 ;
        RECT 68.290 22.495 68.520 24.015 ;
        RECT 68.765 23.005 68.955 24.105 ;
        RECT 69.720 24.005 69.990 24.105 ;
        RECT 69.760 23.975 69.950 24.005 ;
        RECT 86.630 23.950 87.090 24.180 ;
        RECT 102.225 24.295 102.495 24.385 ;
        RECT 103.260 24.295 103.450 25.390 ;
        RECT 102.225 24.105 103.450 24.295 ;
        RECT 102.225 24.005 102.495 24.105 ;
        RECT 102.265 23.975 102.455 24.005 ;
        RECT 86.260 23.140 86.580 23.790 ;
        RECT 69.720 23.005 69.990 23.095 ;
        RECT 68.765 22.815 69.990 23.005 ;
        RECT 86.745 22.980 86.975 23.950 ;
        RECT 87.140 23.140 87.460 23.790 ;
        RECT 68.765 22.765 68.990 22.815 ;
        RECT 67.660 22.095 68.520 22.495 ;
        RECT 68.730 22.445 68.990 22.765 ;
        RECT 69.720 22.715 69.990 22.815 ;
        RECT 86.630 22.750 87.090 22.980 ;
        RECT 69.760 22.685 69.950 22.715 ;
        RECT 87.230 22.545 87.460 23.140 ;
        RECT 102.225 23.005 102.495 23.095 ;
        RECT 103.260 23.005 103.450 24.105 ;
        RECT 103.600 25.185 104.555 25.590 ;
        RECT 104.985 25.590 105.215 27.345 ;
        RECT 105.575 27.335 105.805 27.345 ;
        RECT 105.385 26.735 105.985 27.335 ;
        RECT 104.985 25.345 105.310 25.590 ;
        RECT 105.575 25.585 105.805 26.735 ;
        RECT 103.600 24.415 104.955 25.185 ;
        RECT 103.600 24.025 104.555 24.415 ;
        RECT 105.120 24.255 105.310 25.345 ;
        RECT 103.600 24.015 103.925 24.025 ;
        RECT 102.225 22.815 103.450 23.005 ;
        RECT 102.225 22.715 102.495 22.815 ;
        RECT 103.225 22.765 103.450 22.815 ;
        RECT 102.265 22.685 102.455 22.715 ;
        RECT 86.170 22.255 87.550 22.545 ;
        RECT 103.225 22.445 103.485 22.765 ;
        RECT 103.695 22.495 103.925 24.015 ;
        RECT 104.360 22.495 104.555 24.025 ;
        RECT 104.985 24.000 105.310 24.255 ;
        RECT 105.490 25.345 105.805 25.585 ;
        RECT 105.490 24.255 105.680 25.345 ;
        RECT 106.240 25.185 106.430 27.505 ;
        RECT 106.865 25.585 107.095 27.345 ;
        RECT 107.455 27.335 107.685 27.345 ;
        RECT 107.265 26.735 107.865 27.335 ;
        RECT 107.455 25.590 107.685 26.735 ;
        RECT 106.865 25.345 107.190 25.585 ;
        RECT 105.835 24.415 106.835 25.185 ;
        RECT 105.490 24.000 105.805 24.255 ;
        RECT 104.985 22.855 105.215 24.000 ;
        RECT 56.000 21.865 56.960 22.095 ;
        RECT 57.880 21.890 59.100 22.095 ;
        RECT 57.880 21.865 58.840 21.890 ;
        RECT 59.760 21.865 60.720 22.095 ;
        RECT 61.640 21.865 62.600 22.095 ;
        RECT 56.030 21.815 56.930 21.865 ;
        RECT 57.910 21.815 58.810 21.865 ;
        RECT 63.500 21.775 64.500 22.095 ;
        RECT 65.380 21.775 66.380 22.095 ;
        RECT 67.260 21.865 68.520 22.095 ;
        RECT 103.695 22.095 104.555 22.495 ;
        RECT 104.695 22.255 105.295 22.855 ;
        RECT 105.575 22.255 105.805 24.000 ;
        RECT 106.240 22.095 106.430 24.415 ;
        RECT 107.000 24.255 107.190 25.345 ;
        RECT 106.865 24.000 107.190 24.255 ;
        RECT 107.370 25.345 107.685 25.590 ;
        RECT 107.370 24.255 107.560 25.345 ;
        RECT 108.120 25.185 108.310 27.505 ;
        RECT 109.240 27.345 109.430 28.055 ;
        RECT 109.615 27.505 110.575 27.735 ;
        RECT 111.495 27.505 112.455 27.735 ;
        RECT 108.745 25.585 108.975 27.345 ;
        RECT 109.240 27.100 109.565 27.345 ;
        RECT 109.335 25.590 109.565 27.100 ;
        RECT 108.745 25.345 109.060 25.585 ;
        RECT 107.715 24.415 108.715 25.185 ;
        RECT 107.370 24.010 107.685 24.255 ;
        RECT 106.865 22.855 107.095 24.000 ;
        RECT 106.575 22.255 107.175 22.855 ;
        RECT 107.455 22.255 107.685 24.010 ;
        RECT 108.120 22.095 108.310 24.415 ;
        RECT 108.870 24.255 109.060 25.345 ;
        RECT 108.745 24.010 109.060 24.255 ;
        RECT 109.250 25.345 109.565 25.590 ;
        RECT 109.250 24.255 109.440 25.345 ;
        RECT 110.000 25.185 110.190 27.505 ;
        RECT 110.625 27.295 110.855 27.345 ;
        RECT 111.215 27.295 111.445 27.345 ;
        RECT 110.625 27.105 111.445 27.295 ;
        RECT 110.625 25.585 110.855 27.105 ;
        RECT 111.215 25.585 111.445 27.105 ;
        RECT 110.625 25.345 111.445 25.585 ;
        RECT 109.615 24.415 110.575 25.185 ;
        RECT 109.250 24.015 109.565 24.255 ;
        RECT 108.745 22.855 108.975 24.010 ;
        RECT 108.455 22.255 109.055 22.855 ;
        RECT 109.335 22.255 109.565 24.015 ;
        RECT 110.000 22.095 110.190 24.415 ;
        RECT 110.750 24.255 111.310 25.345 ;
        RECT 111.880 25.185 112.070 27.505 ;
        RECT 112.645 27.345 112.835 28.495 ;
        RECT 112.505 27.335 112.835 27.345 ;
        RECT 112.225 26.735 112.835 27.335 ;
        RECT 113.010 28.495 113.325 28.740 ;
        RECT 113.010 27.735 113.200 28.495 ;
        RECT 113.760 28.290 113.950 32.700 ;
        RECT 114.510 32.495 115.050 32.985 ;
        RECT 115.315 32.930 116.155 33.240 ;
        RECT 115.255 32.700 116.215 32.930 ;
        RECT 114.385 32.255 115.205 32.495 ;
        RECT 114.385 28.735 114.615 32.255 ;
        RECT 114.860 32.250 115.205 32.255 ;
        RECT 114.975 28.735 115.205 32.250 ;
        RECT 114.385 28.545 115.205 28.735 ;
        RECT 114.385 28.495 114.615 28.545 ;
        RECT 114.975 28.495 115.205 28.545 ;
        RECT 115.640 28.290 115.830 32.700 ;
        RECT 116.390 32.495 116.580 33.675 ;
        RECT 116.265 32.250 116.580 32.495 ;
        RECT 116.265 29.095 116.495 32.250 ;
        RECT 116.035 28.495 116.635 29.095 ;
        RECT 113.375 28.060 114.335 28.290 ;
        RECT 115.255 28.060 116.215 28.290 ;
        RECT 113.010 27.715 114.335 27.735 ;
        RECT 115.255 27.715 116.215 27.735 ;
        RECT 113.010 27.525 116.215 27.715 ;
        RECT 113.010 27.505 114.335 27.525 ;
        RECT 115.255 27.505 116.215 27.525 ;
        RECT 113.010 27.100 113.955 27.505 ;
        RECT 113.015 27.095 113.955 27.100 ;
        RECT 114.385 27.295 114.615 27.345 ;
        RECT 114.975 27.295 115.205 27.345 ;
        RECT 114.385 27.105 115.205 27.295 ;
        RECT 112.505 25.585 112.735 26.735 ;
        RECT 113.095 25.585 113.325 27.095 ;
        RECT 113.760 25.585 113.950 27.095 ;
        RECT 112.505 25.345 112.820 25.585 ;
        RECT 111.495 24.415 112.455 25.185 ;
        RECT 110.625 24.015 111.445 24.255 ;
        RECT 110.625 22.495 110.855 24.015 ;
        RECT 111.215 22.495 111.445 24.015 ;
        RECT 110.625 22.305 111.445 22.495 ;
        RECT 110.625 22.255 110.855 22.305 ;
        RECT 111.215 22.255 111.445 22.305 ;
        RECT 111.880 22.095 112.070 24.415 ;
        RECT 112.630 24.255 112.820 25.345 ;
        RECT 112.505 24.000 112.820 24.255 ;
        RECT 113.000 25.195 113.950 25.585 ;
        RECT 114.385 25.585 114.615 27.105 ;
        RECT 114.975 25.585 115.205 27.105 ;
        RECT 114.385 25.345 115.205 25.585 ;
        RECT 113.000 24.415 114.335 25.195 ;
        RECT 113.000 24.015 113.950 24.415 ;
        RECT 114.520 24.255 115.085 25.345 ;
        RECT 115.640 25.185 115.830 27.505 ;
        RECT 116.440 27.345 116.635 28.495 ;
        RECT 116.035 26.735 116.635 27.345 ;
        RECT 116.265 25.585 116.495 26.735 ;
        RECT 116.265 25.345 116.580 25.585 ;
        RECT 115.255 24.415 116.215 25.185 ;
        RECT 113.000 24.010 113.325 24.015 ;
        RECT 112.505 22.255 112.735 24.000 ;
        RECT 113.095 22.485 113.325 24.010 ;
        RECT 113.760 22.485 113.950 24.015 ;
        RECT 114.385 24.005 115.205 24.255 ;
        RECT 114.385 22.885 114.615 24.005 ;
        RECT 114.975 22.885 115.205 24.005 ;
        RECT 113.095 22.255 113.955 22.485 ;
        RECT 114.385 22.285 115.205 22.885 ;
        RECT 114.385 22.255 114.615 22.285 ;
        RECT 114.975 22.255 115.205 22.285 ;
        RECT 113.115 22.135 113.955 22.255 ;
        RECT 115.640 22.135 115.830 24.415 ;
        RECT 116.390 24.255 116.580 25.345 ;
        RECT 116.265 24.020 116.580 24.255 ;
        RECT 116.265 22.255 116.495 24.020 ;
        RECT 113.115 22.095 114.305 22.135 ;
        RECT 115.285 22.095 116.185 22.135 ;
        RECT 103.695 21.865 104.955 22.095 ;
        RECT 67.260 21.775 68.260 21.865 ;
        RECT 103.955 21.775 104.955 21.865 ;
        RECT 105.835 21.775 106.835 22.095 ;
        RECT 107.715 21.775 108.715 22.095 ;
        RECT 109.615 21.865 110.575 22.095 ;
        RECT 111.495 21.865 112.455 22.095 ;
        RECT 113.115 21.890 114.335 22.095 ;
        RECT 113.375 21.865 114.335 21.890 ;
        RECT 115.255 21.865 116.215 22.095 ;
        RECT 113.405 21.815 114.305 21.865 ;
        RECT 115.285 21.815 116.185 21.865 ;
        RECT 0.000 0.000 1.000 1.000 ;
        RECT 144.360 0.000 145.360 1.000 ;
      LAYER met2 ;
        RECT 15.005 223.370 15.355 223.395 ;
        RECT 17.765 223.370 18.115 223.395 ;
        RECT 20.525 223.370 20.875 223.395 ;
        RECT 23.285 223.370 23.635 223.395 ;
        RECT 26.045 223.370 26.395 223.395 ;
        RECT 28.805 223.370 29.155 223.395 ;
        RECT 31.565 223.370 31.915 223.395 ;
        RECT 34.325 223.370 34.675 223.395 ;
        RECT 37.085 223.370 37.435 223.395 ;
        RECT 39.845 223.370 40.195 223.395 ;
        RECT 42.605 223.370 42.955 223.395 ;
        RECT 45.365 223.370 45.715 223.395 ;
        RECT 48.125 223.370 48.475 223.395 ;
        RECT 50.885 223.370 51.235 223.395 ;
        RECT 53.645 223.370 53.995 223.395 ;
        RECT 56.405 223.370 56.755 223.395 ;
        RECT 59.165 223.370 59.515 223.395 ;
        RECT 61.925 223.370 62.275 223.395 ;
        RECT 64.685 223.370 65.035 223.395 ;
        RECT 67.445 223.370 67.795 223.395 ;
        RECT 70.205 223.370 70.555 223.395 ;
        RECT 72.965 223.370 73.315 223.395 ;
        RECT 75.725 223.370 76.075 223.395 ;
        RECT 78.485 223.370 78.835 223.395 ;
        RECT 103.325 223.370 103.675 223.395 ;
        RECT 106.085 223.370 106.435 223.395 ;
        RECT 108.845 223.370 109.195 223.395 ;
        RECT 111.605 223.370 111.955 223.395 ;
        RECT 114.365 223.370 114.715 223.395 ;
        RECT 117.125 223.370 117.475 223.395 ;
        RECT 119.885 223.370 120.235 223.395 ;
        RECT 122.645 223.370 122.995 223.395 ;
        RECT 14.985 223.070 15.375 223.370 ;
        RECT 17.745 223.070 18.135 223.370 ;
        RECT 20.505 223.070 20.895 223.370 ;
        RECT 23.265 223.070 23.655 223.370 ;
        RECT 26.025 223.070 26.415 223.370 ;
        RECT 28.785 223.070 29.175 223.370 ;
        RECT 31.545 223.070 31.935 223.370 ;
        RECT 34.305 223.070 34.695 223.370 ;
        RECT 37.065 223.070 37.455 223.370 ;
        RECT 39.825 223.070 40.215 223.370 ;
        RECT 42.585 223.070 42.975 223.370 ;
        RECT 45.345 223.070 45.735 223.370 ;
        RECT 48.105 223.070 48.495 223.370 ;
        RECT 50.865 223.070 51.255 223.370 ;
        RECT 53.625 223.070 54.015 223.370 ;
        RECT 56.385 223.070 56.775 223.370 ;
        RECT 59.145 223.070 59.535 223.370 ;
        RECT 61.905 223.070 62.295 223.370 ;
        RECT 64.665 223.070 65.055 223.370 ;
        RECT 67.425 223.070 67.815 223.370 ;
        RECT 70.185 223.070 70.575 223.370 ;
        RECT 72.945 223.070 73.335 223.370 ;
        RECT 75.705 223.070 76.095 223.370 ;
        RECT 78.465 223.070 78.855 223.370 ;
        RECT 103.305 223.070 103.695 223.370 ;
        RECT 106.065 223.070 106.455 223.370 ;
        RECT 108.825 223.070 109.215 223.370 ;
        RECT 111.585 223.070 111.975 223.370 ;
        RECT 114.345 223.070 114.735 223.370 ;
        RECT 117.105 223.070 117.495 223.370 ;
        RECT 119.865 223.070 120.255 223.370 ;
        RECT 122.625 223.070 123.015 223.370 ;
        RECT 15.005 220.410 15.355 223.070 ;
        RECT 15.000 218.705 15.355 220.410 ;
        RECT 14.200 218.355 15.355 218.705 ;
        RECT 13.320 206.710 13.620 206.755 ;
        RECT 13.290 206.410 13.650 206.710 ;
        RECT 13.320 206.365 13.620 206.410 ;
        RECT 14.200 205.470 14.550 218.355 ;
        RECT 17.765 217.705 18.115 223.070 ;
        RECT 15.700 217.355 18.115 217.705 ;
        RECT 14.820 206.710 15.120 206.755 ;
        RECT 14.790 206.410 15.150 206.710 ;
        RECT 14.820 206.365 15.120 206.410 ;
        RECT 15.700 205.470 16.050 217.355 ;
        RECT 20.525 216.705 20.875 223.070 ;
        RECT 17.200 216.355 20.875 216.705 ;
        RECT 16.320 206.710 16.620 206.755 ;
        RECT 16.290 206.410 16.650 206.710 ;
        RECT 16.320 206.365 16.620 206.410 ;
        RECT 17.200 205.470 17.550 216.355 ;
        RECT 23.285 215.705 23.635 223.070 ;
        RECT 18.700 215.355 23.635 215.705 ;
        RECT 17.820 206.710 18.120 206.755 ;
        RECT 17.790 206.410 18.150 206.710 ;
        RECT 17.820 206.365 18.120 206.410 ;
        RECT 18.700 205.470 19.050 215.355 ;
        RECT 26.045 214.705 26.395 223.070 ;
        RECT 20.200 214.355 26.395 214.705 ;
        RECT 19.320 206.710 19.620 206.755 ;
        RECT 19.290 206.410 19.650 206.710 ;
        RECT 19.320 206.365 19.620 206.410 ;
        RECT 20.200 205.470 20.550 214.355 ;
        RECT 28.805 213.705 29.155 223.070 ;
        RECT 21.700 213.355 29.155 213.705 ;
        RECT 20.820 206.710 21.120 206.755 ;
        RECT 20.790 206.410 21.150 206.710 ;
        RECT 20.820 206.365 21.120 206.410 ;
        RECT 21.700 205.470 22.050 213.355 ;
        RECT 31.565 212.705 31.915 223.070 ;
        RECT 23.200 212.355 31.915 212.705 ;
        RECT 22.320 206.710 22.620 206.755 ;
        RECT 22.290 206.410 22.650 206.710 ;
        RECT 22.320 206.365 22.620 206.410 ;
        RECT 23.200 205.470 23.550 212.355 ;
        RECT 34.325 211.705 34.675 223.070 ;
        RECT 24.700 211.355 34.675 211.705 ;
        RECT 37.085 211.705 37.435 223.070 ;
        RECT 39.845 212.705 40.195 223.070 ;
        RECT 42.605 216.705 42.955 223.070 ;
        RECT 42.290 216.355 42.955 216.705 ;
        RECT 39.845 212.365 41.140 212.705 ;
        RECT 40.040 212.355 41.140 212.365 ;
        RECT 37.085 211.355 39.640 211.705 ;
        RECT 23.820 206.710 24.120 206.755 ;
        RECT 23.790 206.410 24.150 206.710 ;
        RECT 23.820 206.365 24.120 206.410 ;
        RECT 24.700 205.470 25.050 211.355 ;
        RECT 38.605 208.130 38.905 208.180 ;
        RECT 38.580 207.840 38.930 208.130 ;
        RECT 38.605 207.790 38.905 207.840 ;
        RECT 39.290 206.925 39.640 211.355 ;
        RECT 40.230 208.115 40.530 208.180 ;
        RECT 40.220 207.855 40.540 208.115 ;
        RECT 40.230 207.790 40.530 207.855 ;
        RECT 40.790 206.925 41.140 212.355 ;
        RECT 41.730 208.115 42.030 208.180 ;
        RECT 41.720 207.855 42.040 208.115 ;
        RECT 41.730 207.790 42.030 207.855 ;
        RECT 42.290 206.925 42.640 216.355 ;
        RECT 45.365 215.705 45.715 223.070 ;
        RECT 43.790 215.355 45.715 215.705 ;
        RECT 43.230 208.115 43.530 208.180 ;
        RECT 43.220 207.855 43.540 208.115 ;
        RECT 43.230 207.790 43.530 207.855 ;
        RECT 43.790 206.925 44.140 215.355 ;
        RECT 48.125 214.705 48.475 223.070 ;
        RECT 45.290 214.355 48.475 214.705 ;
        RECT 44.730 208.115 45.030 208.180 ;
        RECT 44.720 207.855 45.040 208.115 ;
        RECT 44.730 207.790 45.030 207.855 ;
        RECT 45.290 206.925 45.640 214.355 ;
        RECT 50.885 213.705 51.235 223.070 ;
        RECT 46.790 213.355 51.235 213.705 ;
        RECT 46.230 208.115 46.530 208.180 ;
        RECT 46.220 207.855 46.540 208.115 ;
        RECT 46.230 207.790 46.530 207.855 ;
        RECT 46.790 206.925 47.140 213.355 ;
        RECT 53.645 212.705 53.995 223.070 ;
        RECT 48.290 212.355 53.995 212.705 ;
        RECT 47.730 208.115 48.030 208.180 ;
        RECT 47.720 207.855 48.040 208.115 ;
        RECT 47.730 207.790 48.030 207.855 ;
        RECT 48.290 206.925 48.640 212.355 ;
        RECT 56.405 211.705 56.755 223.070 ;
        RECT 49.790 211.355 56.755 211.705 ;
        RECT 59.165 211.705 59.515 223.070 ;
        RECT 61.925 212.705 62.275 223.070 ;
        RECT 64.685 213.705 65.035 223.070 ;
        RECT 67.445 214.705 67.795 223.070 ;
        RECT 70.205 215.705 70.555 223.070 ;
        RECT 70.205 215.355 71.640 215.705 ;
        RECT 67.445 214.355 70.140 214.705 ;
        RECT 64.685 213.355 68.640 213.705 ;
        RECT 61.925 212.355 67.140 212.705 ;
        RECT 59.165 211.355 65.640 211.705 ;
        RECT 49.230 208.115 49.530 208.180 ;
        RECT 49.220 207.855 49.540 208.115 ;
        RECT 49.230 207.790 49.530 207.855 ;
        RECT 49.790 206.925 50.140 211.355 ;
        RECT 50.730 208.115 51.030 208.180 ;
        RECT 51.385 208.130 51.685 208.180 ;
        RECT 64.605 208.130 64.905 208.180 ;
        RECT 50.720 207.855 51.040 208.115 ;
        RECT 50.730 207.790 51.030 207.855 ;
        RECT 51.360 207.840 51.710 208.130 ;
        RECT 64.580 207.840 64.930 208.130 ;
        RECT 51.385 207.790 51.685 207.840 ;
        RECT 64.605 207.790 64.905 207.840 ;
        RECT 65.290 206.925 65.640 211.355 ;
        RECT 66.230 208.115 66.530 208.180 ;
        RECT 66.220 207.855 66.540 208.115 ;
        RECT 66.230 207.790 66.530 207.855 ;
        RECT 66.790 206.925 67.140 212.355 ;
        RECT 67.730 208.115 68.030 208.180 ;
        RECT 67.720 207.855 68.040 208.115 ;
        RECT 67.730 207.790 68.030 207.855 ;
        RECT 68.290 206.925 68.640 213.355 ;
        RECT 69.230 208.115 69.530 208.180 ;
        RECT 69.220 207.855 69.540 208.115 ;
        RECT 69.230 207.790 69.530 207.855 ;
        RECT 69.790 206.925 70.140 214.355 ;
        RECT 70.730 208.115 71.030 208.180 ;
        RECT 70.720 207.855 71.040 208.115 ;
        RECT 70.730 207.790 71.030 207.855 ;
        RECT 71.290 206.925 71.640 215.355 ;
        RECT 72.965 213.705 73.315 223.070 ;
        RECT 72.790 213.355 73.315 213.705 ;
        RECT 72.230 208.115 72.530 208.180 ;
        RECT 72.220 207.855 72.540 208.115 ;
        RECT 72.230 207.790 72.530 207.855 ;
        RECT 72.790 206.925 73.140 213.355 ;
        RECT 75.725 212.705 76.075 223.070 ;
        RECT 74.290 212.355 76.075 212.705 ;
        RECT 73.730 208.115 74.030 208.180 ;
        RECT 73.720 207.855 74.040 208.115 ;
        RECT 73.730 207.790 74.030 207.855 ;
        RECT 74.290 206.925 74.640 212.355 ;
        RECT 75.790 211.700 76.140 211.705 ;
        RECT 78.485 211.700 78.835 223.070 ;
        RECT 75.790 211.355 78.835 211.700 ;
        RECT 103.325 211.705 103.675 223.070 ;
        RECT 106.085 212.705 106.435 223.070 ;
        RECT 108.845 213.705 109.195 223.070 ;
        RECT 111.605 214.705 111.955 223.070 ;
        RECT 114.365 214.705 114.715 223.070 ;
        RECT 111.605 214.355 112.595 214.705 ;
        RECT 108.845 213.355 111.095 213.705 ;
        RECT 106.085 212.355 109.595 212.705 ;
        RECT 103.325 211.355 108.095 211.705 ;
        RECT 75.790 211.350 78.640 211.355 ;
        RECT 75.230 208.115 75.530 208.180 ;
        RECT 75.220 207.855 75.540 208.115 ;
        RECT 75.230 207.790 75.530 207.855 ;
        RECT 75.790 206.925 76.140 211.350 ;
        RECT 76.730 208.115 77.030 208.180 ;
        RECT 77.385 208.130 77.685 208.180 ;
        RECT 76.720 207.855 77.040 208.115 ;
        RECT 76.730 207.790 77.030 207.855 ;
        RECT 77.360 207.840 77.710 208.130 ;
        RECT 77.385 207.790 77.685 207.840 ;
        RECT 106.755 206.625 107.055 206.675 ;
        RECT 39.760 206.190 40.080 206.450 ;
        RECT 41.260 206.190 41.580 206.450 ;
        RECT 42.760 206.190 43.080 206.450 ;
        RECT 44.260 206.190 44.580 206.450 ;
        RECT 45.760 206.190 46.080 206.450 ;
        RECT 47.260 206.190 47.580 206.450 ;
        RECT 48.760 206.190 49.080 206.450 ;
        RECT 50.260 206.190 50.580 206.450 ;
        RECT 65.760 206.190 66.080 206.450 ;
        RECT 67.260 206.190 67.580 206.450 ;
        RECT 68.760 206.190 69.080 206.450 ;
        RECT 70.260 206.190 70.580 206.450 ;
        RECT 71.760 206.190 72.080 206.450 ;
        RECT 73.260 206.190 73.580 206.450 ;
        RECT 74.760 206.190 75.080 206.450 ;
        RECT 76.260 206.190 76.580 206.450 ;
        RECT 106.730 206.335 107.080 206.625 ;
        RECT 107.245 206.610 107.545 206.675 ;
        RECT 107.235 206.350 107.555 206.610 ;
        RECT 106.755 206.285 107.055 206.335 ;
        RECT 107.245 206.285 107.545 206.350 ;
        RECT 39.835 205.505 40.005 206.190 ;
        RECT 41.335 205.505 41.505 206.190 ;
        RECT 42.835 205.505 43.005 206.190 ;
        RECT 44.335 205.505 44.505 206.190 ;
        RECT 45.835 205.505 46.005 206.190 ;
        RECT 47.335 205.505 47.505 206.190 ;
        RECT 48.835 205.505 49.005 206.190 ;
        RECT 50.335 205.505 50.505 206.190 ;
        RECT 65.835 205.505 66.005 206.190 ;
        RECT 67.335 205.505 67.505 206.190 ;
        RECT 68.835 205.505 69.005 206.190 ;
        RECT 70.335 205.505 70.505 206.190 ;
        RECT 71.835 205.505 72.005 206.190 ;
        RECT 73.335 205.505 73.505 206.190 ;
        RECT 74.835 205.505 75.005 206.190 ;
        RECT 76.335 205.505 76.505 206.190 ;
        RECT 107.745 206.135 108.095 211.355 ;
        RECT 108.745 206.610 109.045 206.675 ;
        RECT 108.735 206.350 109.055 206.610 ;
        RECT 108.745 206.285 109.045 206.350 ;
        RECT 109.245 206.135 109.595 212.355 ;
        RECT 110.245 206.610 110.545 206.675 ;
        RECT 110.235 206.350 110.555 206.610 ;
        RECT 110.245 206.285 110.545 206.350 ;
        RECT 110.745 206.135 111.095 213.355 ;
        RECT 111.745 206.610 112.045 206.675 ;
        RECT 111.735 206.350 112.055 206.610 ;
        RECT 111.745 206.285 112.045 206.350 ;
        RECT 112.245 206.135 112.595 214.355 ;
        RECT 113.745 214.355 114.715 214.705 ;
        RECT 113.245 206.610 113.545 206.675 ;
        RECT 113.235 206.350 113.555 206.610 ;
        RECT 113.245 206.285 113.545 206.350 ;
        RECT 113.745 206.135 114.095 214.355 ;
        RECT 117.125 213.705 117.475 223.070 ;
        RECT 115.245 213.355 117.475 213.705 ;
        RECT 114.745 206.610 115.045 206.675 ;
        RECT 114.735 206.350 115.055 206.610 ;
        RECT 114.745 206.285 115.045 206.350 ;
        RECT 115.245 206.135 115.595 213.355 ;
        RECT 119.885 212.705 120.235 223.070 ;
        RECT 116.745 212.355 120.235 212.705 ;
        RECT 116.245 206.610 116.545 206.675 ;
        RECT 116.235 206.350 116.555 206.610 ;
        RECT 116.245 206.285 116.545 206.350 ;
        RECT 116.745 206.135 117.095 212.355 ;
        RECT 122.645 211.705 122.995 223.070 ;
        RECT 118.245 211.355 122.995 211.705 ;
        RECT 117.745 206.610 118.045 206.675 ;
        RECT 117.735 206.350 118.055 206.610 ;
        RECT 117.745 206.285 118.045 206.350 ;
        RECT 118.245 206.135 118.595 211.355 ;
        RECT 119.285 206.625 119.585 206.675 ;
        RECT 119.260 206.335 119.610 206.625 ;
        RECT 119.285 206.285 119.585 206.335 ;
        RECT 107.720 205.735 108.120 206.135 ;
        RECT 109.220 205.735 109.620 206.135 ;
        RECT 110.720 205.735 111.120 206.135 ;
        RECT 112.220 205.735 112.620 206.135 ;
        RECT 113.720 205.735 114.120 206.135 ;
        RECT 115.220 205.735 115.620 206.135 ;
        RECT 116.720 205.735 117.120 206.135 ;
        RECT 118.220 205.735 118.620 206.135 ;
        RECT 39.835 205.335 40.460 205.505 ;
        RECT 41.335 205.335 41.960 205.505 ;
        RECT 42.835 205.335 43.460 205.505 ;
        RECT 44.335 205.335 44.960 205.505 ;
        RECT 45.835 205.335 46.460 205.505 ;
        RECT 47.335 205.335 47.960 205.505 ;
        RECT 48.835 205.335 49.460 205.505 ;
        RECT 50.335 205.335 50.960 205.505 ;
        RECT 65.835 205.335 66.460 205.505 ;
        RECT 67.335 205.335 67.960 205.505 ;
        RECT 68.835 205.335 69.460 205.505 ;
        RECT 70.335 205.335 70.960 205.505 ;
        RECT 71.835 205.335 72.460 205.505 ;
        RECT 73.335 205.335 73.960 205.505 ;
        RECT 74.835 205.335 75.460 205.505 ;
        RECT 76.335 205.335 76.960 205.505 ;
        RECT 39.335 203.315 39.595 203.390 ;
        RECT 39.335 203.145 40.005 203.315 ;
        RECT 39.335 203.070 39.595 203.145 ;
        RECT 39.240 202.830 39.500 202.905 ;
        RECT 39.240 202.585 39.550 202.830 ;
        RECT 38.725 202.500 39.075 202.545 ;
        RECT 38.695 202.150 39.105 202.500 ;
        RECT 38.725 202.105 39.075 202.150 ;
        RECT 38.580 201.450 38.930 201.495 ;
        RECT 38.550 201.100 38.960 201.450 ;
        RECT 13.315 201.030 13.615 201.095 ;
        RECT 14.815 201.030 15.115 201.095 ;
        RECT 16.315 201.030 16.615 201.095 ;
        RECT 17.815 201.030 18.115 201.095 ;
        RECT 19.315 201.030 19.615 201.095 ;
        RECT 20.815 201.030 21.115 201.095 ;
        RECT 22.315 201.030 22.615 201.095 ;
        RECT 23.815 201.030 24.115 201.095 ;
        RECT 38.580 201.055 38.930 201.100 ;
        RECT 13.305 200.770 13.625 201.030 ;
        RECT 14.805 200.770 15.125 201.030 ;
        RECT 16.305 200.770 16.625 201.030 ;
        RECT 17.805 200.770 18.125 201.030 ;
        RECT 19.305 200.770 19.625 201.030 ;
        RECT 20.805 200.770 21.125 201.030 ;
        RECT 22.305 200.770 22.625 201.030 ;
        RECT 23.805 200.770 24.125 201.030 ;
        RECT 13.315 200.705 13.615 200.770 ;
        RECT 14.815 200.705 15.115 200.770 ;
        RECT 16.315 200.705 16.615 200.770 ;
        RECT 17.815 200.705 18.115 200.770 ;
        RECT 19.315 200.705 19.615 200.770 ;
        RECT 20.815 200.705 21.115 200.770 ;
        RECT 22.315 200.705 22.615 200.770 ;
        RECT 23.815 200.705 24.115 200.770 ;
        RECT 39.380 200.520 39.550 202.585 ;
        RECT 39.305 200.260 39.625 200.520 ;
        RECT 39.835 199.365 40.005 203.145 ;
        RECT 39.790 199.045 40.050 199.365 ;
        RECT 40.290 198.835 40.460 205.335 ;
        RECT 40.835 203.315 41.095 203.390 ;
        RECT 40.835 203.145 41.505 203.315 ;
        RECT 40.835 203.070 41.095 203.145 ;
        RECT 40.740 202.830 41.000 202.905 ;
        RECT 40.740 202.585 41.050 202.830 ;
        RECT 40.880 200.520 41.050 202.585 ;
        RECT 40.805 200.260 41.125 200.520 ;
        RECT 41.335 199.365 41.505 203.145 ;
        RECT 41.290 199.045 41.550 199.365 ;
        RECT 41.790 198.835 41.960 205.335 ;
        RECT 42.335 203.315 42.595 203.390 ;
        RECT 42.335 203.145 43.005 203.315 ;
        RECT 42.335 203.070 42.595 203.145 ;
        RECT 42.240 202.830 42.500 202.905 ;
        RECT 42.240 202.585 42.550 202.830 ;
        RECT 42.380 200.520 42.550 202.585 ;
        RECT 42.305 200.260 42.625 200.520 ;
        RECT 42.835 199.365 43.005 203.145 ;
        RECT 42.790 199.045 43.050 199.365 ;
        RECT 43.290 198.835 43.460 205.335 ;
        RECT 43.835 203.315 44.095 203.390 ;
        RECT 43.835 203.145 44.505 203.315 ;
        RECT 43.835 203.070 44.095 203.145 ;
        RECT 43.740 202.830 44.000 202.905 ;
        RECT 43.740 202.585 44.050 202.830 ;
        RECT 43.880 200.520 44.050 202.585 ;
        RECT 43.805 200.260 44.125 200.520 ;
        RECT 44.335 199.365 44.505 203.145 ;
        RECT 44.290 199.045 44.550 199.365 ;
        RECT 44.790 198.835 44.960 205.335 ;
        RECT 45.335 203.315 45.595 203.390 ;
        RECT 45.335 203.145 46.005 203.315 ;
        RECT 45.335 203.070 45.595 203.145 ;
        RECT 45.240 202.830 45.500 202.905 ;
        RECT 45.240 202.585 45.550 202.830 ;
        RECT 45.380 200.520 45.550 202.585 ;
        RECT 45.305 200.260 45.625 200.520 ;
        RECT 45.835 199.365 46.005 203.145 ;
        RECT 45.790 199.045 46.050 199.365 ;
        RECT 46.290 198.835 46.460 205.335 ;
        RECT 46.835 203.315 47.095 203.390 ;
        RECT 46.835 203.145 47.505 203.315 ;
        RECT 46.835 203.070 47.095 203.145 ;
        RECT 46.740 202.830 47.000 202.905 ;
        RECT 46.740 202.585 47.050 202.830 ;
        RECT 46.880 200.520 47.050 202.585 ;
        RECT 46.805 200.260 47.125 200.520 ;
        RECT 47.335 199.365 47.505 203.145 ;
        RECT 47.290 199.045 47.550 199.365 ;
        RECT 47.790 198.835 47.960 205.335 ;
        RECT 48.335 203.315 48.595 203.390 ;
        RECT 48.335 203.145 49.005 203.315 ;
        RECT 48.335 203.070 48.595 203.145 ;
        RECT 48.240 202.830 48.500 202.905 ;
        RECT 48.240 202.585 48.550 202.830 ;
        RECT 48.380 200.520 48.550 202.585 ;
        RECT 48.305 200.260 48.625 200.520 ;
        RECT 48.835 199.365 49.005 203.145 ;
        RECT 48.790 199.045 49.050 199.365 ;
        RECT 49.290 198.835 49.460 205.335 ;
        RECT 49.835 203.315 50.095 203.390 ;
        RECT 49.835 203.145 50.505 203.315 ;
        RECT 49.835 203.070 50.095 203.145 ;
        RECT 49.740 202.830 50.000 202.905 ;
        RECT 49.740 202.585 50.050 202.830 ;
        RECT 49.880 200.520 50.050 202.585 ;
        RECT 49.805 200.260 50.125 200.520 ;
        RECT 50.335 199.365 50.505 203.145 ;
        RECT 50.290 199.045 50.550 199.365 ;
        RECT 50.790 198.835 50.960 205.335 ;
        RECT 65.335 203.315 65.595 203.390 ;
        RECT 65.335 203.145 66.005 203.315 ;
        RECT 65.335 203.070 65.595 203.145 ;
        RECT 65.240 202.830 65.500 202.905 ;
        RECT 65.240 202.585 65.550 202.830 ;
        RECT 51.260 202.500 51.610 202.545 ;
        RECT 64.725 202.500 65.075 202.545 ;
        RECT 51.230 202.150 51.640 202.500 ;
        RECT 64.695 202.150 65.105 202.500 ;
        RECT 51.260 202.105 51.610 202.150 ;
        RECT 64.725 202.105 65.075 202.150 ;
        RECT 51.360 201.450 51.710 201.495 ;
        RECT 64.580 201.450 64.930 201.495 ;
        RECT 51.330 201.100 51.740 201.450 ;
        RECT 64.550 201.100 64.960 201.450 ;
        RECT 51.360 201.055 51.710 201.100 ;
        RECT 64.580 201.055 64.930 201.100 ;
        RECT 65.380 200.520 65.550 202.585 ;
        RECT 65.305 200.260 65.625 200.520 ;
        RECT 65.835 199.365 66.005 203.145 ;
        RECT 65.790 199.045 66.050 199.365 ;
        RECT 66.290 198.835 66.460 205.335 ;
        RECT 66.835 203.315 67.095 203.390 ;
        RECT 66.835 203.145 67.505 203.315 ;
        RECT 66.835 203.070 67.095 203.145 ;
        RECT 66.740 202.830 67.000 202.905 ;
        RECT 66.740 202.585 67.050 202.830 ;
        RECT 66.880 200.520 67.050 202.585 ;
        RECT 66.805 200.260 67.125 200.520 ;
        RECT 67.335 199.365 67.505 203.145 ;
        RECT 67.290 199.045 67.550 199.365 ;
        RECT 67.790 198.835 67.960 205.335 ;
        RECT 68.335 203.315 68.595 203.390 ;
        RECT 68.335 203.145 69.005 203.315 ;
        RECT 68.335 203.070 68.595 203.145 ;
        RECT 68.240 202.830 68.500 202.905 ;
        RECT 68.240 202.585 68.550 202.830 ;
        RECT 68.380 200.520 68.550 202.585 ;
        RECT 68.305 200.260 68.625 200.520 ;
        RECT 68.835 199.365 69.005 203.145 ;
        RECT 68.790 199.045 69.050 199.365 ;
        RECT 69.290 198.835 69.460 205.335 ;
        RECT 69.835 203.315 70.095 203.390 ;
        RECT 69.835 203.145 70.505 203.315 ;
        RECT 69.835 203.070 70.095 203.145 ;
        RECT 69.740 202.830 70.000 202.905 ;
        RECT 69.740 202.585 70.050 202.830 ;
        RECT 69.880 200.520 70.050 202.585 ;
        RECT 69.805 200.260 70.125 200.520 ;
        RECT 70.335 199.365 70.505 203.145 ;
        RECT 70.290 199.045 70.550 199.365 ;
        RECT 70.790 198.835 70.960 205.335 ;
        RECT 71.335 203.315 71.595 203.390 ;
        RECT 71.335 203.145 72.005 203.315 ;
        RECT 71.335 203.070 71.595 203.145 ;
        RECT 71.240 202.830 71.500 202.905 ;
        RECT 71.240 202.585 71.550 202.830 ;
        RECT 71.380 200.520 71.550 202.585 ;
        RECT 71.305 200.260 71.625 200.520 ;
        RECT 71.835 199.365 72.005 203.145 ;
        RECT 71.790 199.045 72.050 199.365 ;
        RECT 72.290 198.835 72.460 205.335 ;
        RECT 72.835 203.315 73.095 203.390 ;
        RECT 72.835 203.145 73.505 203.315 ;
        RECT 72.835 203.070 73.095 203.145 ;
        RECT 72.740 202.830 73.000 202.905 ;
        RECT 72.740 202.585 73.050 202.830 ;
        RECT 72.880 200.520 73.050 202.585 ;
        RECT 72.805 200.260 73.125 200.520 ;
        RECT 73.335 199.365 73.505 203.145 ;
        RECT 73.290 199.045 73.550 199.365 ;
        RECT 73.790 198.835 73.960 205.335 ;
        RECT 74.335 203.315 74.595 203.390 ;
        RECT 74.335 203.145 75.005 203.315 ;
        RECT 74.335 203.070 74.595 203.145 ;
        RECT 74.240 202.830 74.500 202.905 ;
        RECT 74.240 202.585 74.550 202.830 ;
        RECT 74.380 200.520 74.550 202.585 ;
        RECT 74.305 200.260 74.625 200.520 ;
        RECT 74.835 199.365 75.005 203.145 ;
        RECT 74.790 199.045 75.050 199.365 ;
        RECT 75.290 198.835 75.460 205.335 ;
        RECT 75.835 203.315 76.095 203.390 ;
        RECT 75.835 203.145 76.505 203.315 ;
        RECT 75.835 203.070 76.095 203.145 ;
        RECT 75.740 202.830 76.000 202.905 ;
        RECT 75.740 202.585 76.050 202.830 ;
        RECT 75.880 200.520 76.050 202.585 ;
        RECT 75.805 200.260 76.125 200.520 ;
        RECT 76.335 199.365 76.505 203.145 ;
        RECT 76.290 199.045 76.550 199.365 ;
        RECT 76.790 198.835 76.960 205.335 ;
        RECT 77.260 202.500 77.610 202.545 ;
        RECT 77.230 202.150 77.640 202.500 ;
        RECT 77.260 202.105 77.610 202.150 ;
        RECT 108.245 201.545 108.505 201.865 ;
        RECT 109.745 201.545 110.005 201.865 ;
        RECT 111.245 201.545 111.505 201.865 ;
        RECT 112.745 201.545 113.005 201.865 ;
        RECT 114.245 201.545 114.505 201.865 ;
        RECT 115.745 201.545 116.005 201.865 ;
        RECT 117.245 201.545 117.505 201.865 ;
        RECT 118.745 201.545 119.005 201.865 ;
        RECT 77.360 201.450 77.710 201.495 ;
        RECT 77.330 201.100 77.740 201.450 ;
        RECT 107.790 201.125 108.050 201.445 ;
        RECT 77.360 201.055 77.710 201.100 ;
        RECT 106.655 200.625 106.955 201.015 ;
        RECT 107.315 200.950 107.615 201.015 ;
        RECT 107.305 200.690 107.625 200.950 ;
        RECT 107.315 200.625 107.615 200.690 ;
        RECT 39.380 198.665 40.460 198.835 ;
        RECT 40.880 198.665 41.960 198.835 ;
        RECT 42.380 198.665 43.460 198.835 ;
        RECT 43.880 198.665 44.960 198.835 ;
        RECT 45.380 198.665 46.460 198.835 ;
        RECT 46.880 198.665 47.960 198.835 ;
        RECT 48.380 198.665 49.460 198.835 ;
        RECT 49.880 198.665 50.960 198.835 ;
        RECT 65.380 198.665 66.460 198.835 ;
        RECT 66.880 198.665 67.960 198.835 ;
        RECT 68.380 198.665 69.460 198.835 ;
        RECT 69.880 198.665 70.960 198.835 ;
        RECT 71.380 198.665 72.460 198.835 ;
        RECT 72.880 198.665 73.960 198.835 ;
        RECT 74.380 198.665 75.460 198.835 ;
        RECT 75.880 198.665 76.960 198.835 ;
        RECT 38.755 195.760 39.055 195.810 ;
        RECT 38.730 195.470 39.080 195.760 ;
        RECT 38.755 195.420 39.055 195.470 ;
        RECT 38.605 183.955 38.905 184.005 ;
        RECT 38.580 183.665 38.930 183.955 ;
        RECT 38.605 183.615 38.905 183.665 ;
        RECT 39.380 183.085 39.550 198.665 ;
        RECT 40.215 198.370 40.535 198.415 ;
        RECT 39.835 198.200 40.535 198.370 ;
        RECT 39.835 183.505 40.005 198.200 ;
        RECT 40.215 198.155 40.535 198.200 ;
        RECT 40.225 195.745 40.525 195.810 ;
        RECT 40.215 195.485 40.535 195.745 ;
        RECT 40.225 195.420 40.525 195.485 ;
        RECT 40.225 183.940 40.525 184.005 ;
        RECT 40.215 183.680 40.535 183.940 ;
        RECT 40.225 183.615 40.525 183.680 ;
        RECT 39.790 183.185 40.050 183.505 ;
        RECT 40.880 183.085 41.050 198.665 ;
        RECT 41.715 198.370 42.035 198.415 ;
        RECT 41.335 198.200 42.035 198.370 ;
        RECT 41.335 183.505 41.505 198.200 ;
        RECT 41.715 198.155 42.035 198.200 ;
        RECT 41.725 195.745 42.025 195.810 ;
        RECT 41.715 195.485 42.035 195.745 ;
        RECT 41.725 195.420 42.025 195.485 ;
        RECT 41.725 183.940 42.025 184.005 ;
        RECT 41.715 183.680 42.035 183.940 ;
        RECT 41.725 183.615 42.025 183.680 ;
        RECT 41.290 183.185 41.550 183.505 ;
        RECT 42.380 183.085 42.550 198.665 ;
        RECT 43.215 198.370 43.535 198.415 ;
        RECT 42.835 198.200 43.535 198.370 ;
        RECT 42.835 183.505 43.005 198.200 ;
        RECT 43.215 198.155 43.535 198.200 ;
        RECT 43.225 195.745 43.525 195.810 ;
        RECT 43.215 195.485 43.535 195.745 ;
        RECT 43.225 195.420 43.525 195.485 ;
        RECT 43.225 183.940 43.525 184.005 ;
        RECT 43.215 183.680 43.535 183.940 ;
        RECT 43.225 183.615 43.525 183.680 ;
        RECT 42.790 183.185 43.050 183.505 ;
        RECT 43.880 183.085 44.050 198.665 ;
        RECT 44.715 198.370 45.035 198.415 ;
        RECT 44.335 198.200 45.035 198.370 ;
        RECT 44.335 183.505 44.505 198.200 ;
        RECT 44.715 198.155 45.035 198.200 ;
        RECT 44.725 195.745 45.025 195.810 ;
        RECT 44.715 195.485 45.035 195.745 ;
        RECT 44.725 195.420 45.025 195.485 ;
        RECT 44.725 183.940 45.025 184.005 ;
        RECT 44.715 183.680 45.035 183.940 ;
        RECT 44.725 183.615 45.025 183.680 ;
        RECT 44.290 183.185 44.550 183.505 ;
        RECT 45.380 183.085 45.550 198.665 ;
        RECT 46.215 198.370 46.535 198.415 ;
        RECT 45.835 198.200 46.535 198.370 ;
        RECT 45.835 183.505 46.005 198.200 ;
        RECT 46.215 198.155 46.535 198.200 ;
        RECT 46.225 195.745 46.525 195.810 ;
        RECT 46.215 195.485 46.535 195.745 ;
        RECT 46.225 195.420 46.525 195.485 ;
        RECT 46.225 183.940 46.525 184.005 ;
        RECT 46.215 183.680 46.535 183.940 ;
        RECT 46.225 183.615 46.525 183.680 ;
        RECT 45.790 183.185 46.050 183.505 ;
        RECT 46.880 183.085 47.050 198.665 ;
        RECT 47.715 198.370 48.035 198.415 ;
        RECT 47.335 198.200 48.035 198.370 ;
        RECT 47.335 183.505 47.505 198.200 ;
        RECT 47.715 198.155 48.035 198.200 ;
        RECT 47.725 195.745 48.025 195.810 ;
        RECT 47.715 195.485 48.035 195.745 ;
        RECT 47.725 195.420 48.025 195.485 ;
        RECT 47.725 183.940 48.025 184.005 ;
        RECT 47.715 183.680 48.035 183.940 ;
        RECT 47.725 183.615 48.025 183.680 ;
        RECT 47.290 183.185 47.550 183.505 ;
        RECT 48.380 183.085 48.550 198.665 ;
        RECT 49.215 198.370 49.535 198.415 ;
        RECT 48.835 198.200 49.535 198.370 ;
        RECT 48.835 183.505 49.005 198.200 ;
        RECT 49.215 198.155 49.535 198.200 ;
        RECT 49.225 195.745 49.525 195.810 ;
        RECT 49.215 195.485 49.535 195.745 ;
        RECT 49.225 195.420 49.525 195.485 ;
        RECT 49.225 183.940 49.525 184.005 ;
        RECT 49.215 183.680 49.535 183.940 ;
        RECT 49.225 183.615 49.525 183.680 ;
        RECT 48.790 183.185 49.050 183.505 ;
        RECT 49.880 183.085 50.050 198.665 ;
        RECT 50.715 198.370 51.035 198.415 ;
        RECT 50.335 198.200 51.035 198.370 ;
        RECT 50.335 183.505 50.505 198.200 ;
        RECT 50.715 198.155 51.035 198.200 ;
        RECT 50.725 195.745 51.025 195.810 ;
        RECT 51.285 195.760 51.585 195.810 ;
        RECT 64.755 195.760 65.055 195.810 ;
        RECT 50.715 195.485 51.035 195.745 ;
        RECT 50.725 195.420 51.025 195.485 ;
        RECT 51.260 195.470 51.610 195.760 ;
        RECT 64.730 195.470 65.080 195.760 ;
        RECT 51.285 195.420 51.585 195.470 ;
        RECT 64.755 195.420 65.055 195.470 ;
        RECT 50.725 183.940 51.025 184.005 ;
        RECT 50.715 183.680 51.035 183.940 ;
        RECT 50.725 183.615 51.025 183.680 ;
        RECT 51.385 183.615 51.685 184.005 ;
        RECT 64.605 183.955 64.905 184.005 ;
        RECT 64.580 183.665 64.930 183.955 ;
        RECT 64.605 183.615 64.905 183.665 ;
        RECT 50.290 183.185 50.550 183.505 ;
        RECT 65.380 183.085 65.550 198.665 ;
        RECT 66.215 198.370 66.535 198.415 ;
        RECT 65.835 198.200 66.535 198.370 ;
        RECT 65.835 183.505 66.005 198.200 ;
        RECT 66.215 198.155 66.535 198.200 ;
        RECT 66.225 195.745 66.525 195.810 ;
        RECT 66.215 195.485 66.535 195.745 ;
        RECT 66.225 195.420 66.525 195.485 ;
        RECT 66.225 183.940 66.525 184.005 ;
        RECT 66.215 183.680 66.535 183.940 ;
        RECT 66.225 183.615 66.525 183.680 ;
        RECT 65.790 183.185 66.050 183.505 ;
        RECT 66.880 183.085 67.050 198.665 ;
        RECT 67.715 198.370 68.035 198.415 ;
        RECT 67.335 198.200 68.035 198.370 ;
        RECT 67.335 183.505 67.505 198.200 ;
        RECT 67.715 198.155 68.035 198.200 ;
        RECT 67.725 195.745 68.025 195.810 ;
        RECT 67.715 195.485 68.035 195.745 ;
        RECT 67.725 195.420 68.025 195.485 ;
        RECT 67.725 183.940 68.025 184.005 ;
        RECT 67.715 183.680 68.035 183.940 ;
        RECT 67.725 183.615 68.025 183.680 ;
        RECT 67.290 183.185 67.550 183.505 ;
        RECT 68.380 183.085 68.550 198.665 ;
        RECT 69.215 198.370 69.535 198.415 ;
        RECT 68.835 198.200 69.535 198.370 ;
        RECT 68.835 183.505 69.005 198.200 ;
        RECT 69.215 198.155 69.535 198.200 ;
        RECT 69.225 195.745 69.525 195.810 ;
        RECT 69.215 195.485 69.535 195.745 ;
        RECT 69.225 195.420 69.525 195.485 ;
        RECT 69.225 183.940 69.525 184.005 ;
        RECT 69.215 183.680 69.535 183.940 ;
        RECT 69.225 183.615 69.525 183.680 ;
        RECT 68.790 183.185 69.050 183.505 ;
        RECT 69.880 183.085 70.050 198.665 ;
        RECT 70.715 198.370 71.035 198.415 ;
        RECT 70.335 198.200 71.035 198.370 ;
        RECT 70.335 183.505 70.505 198.200 ;
        RECT 70.715 198.155 71.035 198.200 ;
        RECT 70.725 195.745 71.025 195.810 ;
        RECT 70.715 195.485 71.035 195.745 ;
        RECT 70.725 195.420 71.025 195.485 ;
        RECT 70.725 183.940 71.025 184.005 ;
        RECT 70.715 183.680 71.035 183.940 ;
        RECT 70.725 183.615 71.025 183.680 ;
        RECT 70.290 183.185 70.550 183.505 ;
        RECT 71.380 183.085 71.550 198.665 ;
        RECT 72.215 198.370 72.535 198.415 ;
        RECT 71.835 198.200 72.535 198.370 ;
        RECT 71.835 183.505 72.005 198.200 ;
        RECT 72.215 198.155 72.535 198.200 ;
        RECT 72.225 195.745 72.525 195.810 ;
        RECT 72.215 195.485 72.535 195.745 ;
        RECT 72.225 195.420 72.525 195.485 ;
        RECT 72.225 183.940 72.525 184.005 ;
        RECT 72.215 183.680 72.535 183.940 ;
        RECT 72.225 183.615 72.525 183.680 ;
        RECT 71.790 183.185 72.050 183.505 ;
        RECT 72.880 183.085 73.050 198.665 ;
        RECT 73.715 198.370 74.035 198.415 ;
        RECT 73.335 198.200 74.035 198.370 ;
        RECT 73.335 183.505 73.505 198.200 ;
        RECT 73.715 198.155 74.035 198.200 ;
        RECT 73.725 195.745 74.025 195.810 ;
        RECT 73.715 195.485 74.035 195.745 ;
        RECT 73.725 195.420 74.025 195.485 ;
        RECT 73.725 183.940 74.025 184.005 ;
        RECT 73.715 183.680 74.035 183.940 ;
        RECT 73.725 183.615 74.025 183.680 ;
        RECT 73.290 183.185 73.550 183.505 ;
        RECT 74.380 183.085 74.550 198.665 ;
        RECT 75.215 198.370 75.535 198.415 ;
        RECT 74.835 198.200 75.535 198.370 ;
        RECT 74.835 183.505 75.005 198.200 ;
        RECT 75.215 198.155 75.535 198.200 ;
        RECT 75.225 195.745 75.525 195.810 ;
        RECT 75.215 195.485 75.535 195.745 ;
        RECT 75.225 195.420 75.525 195.485 ;
        RECT 75.225 183.940 75.525 184.005 ;
        RECT 75.215 183.680 75.535 183.940 ;
        RECT 75.225 183.615 75.525 183.680 ;
        RECT 74.790 183.185 75.050 183.505 ;
        RECT 75.880 183.085 76.050 198.665 ;
        RECT 76.715 198.370 77.035 198.415 ;
        RECT 76.335 198.200 77.035 198.370 ;
        RECT 76.335 183.505 76.505 198.200 ;
        RECT 76.715 198.155 77.035 198.200 ;
        RECT 76.725 195.745 77.025 195.810 ;
        RECT 77.285 195.760 77.585 195.810 ;
        RECT 76.715 195.485 77.035 195.745 ;
        RECT 76.725 195.420 77.025 195.485 ;
        RECT 77.260 195.470 77.610 195.760 ;
        RECT 77.285 195.420 77.585 195.470 ;
        RECT 106.755 189.160 107.055 189.210 ;
        RECT 106.730 188.870 107.080 189.160 ;
        RECT 107.315 189.145 107.615 189.210 ;
        RECT 107.305 188.885 107.625 189.145 ;
        RECT 106.755 188.820 107.055 188.870 ;
        RECT 107.315 188.820 107.615 188.885 ;
        RECT 107.305 186.430 107.625 186.475 ;
        RECT 107.835 186.430 108.005 201.125 ;
        RECT 107.305 186.260 108.005 186.430 ;
        RECT 107.305 186.215 107.625 186.260 ;
        RECT 108.290 185.965 108.460 201.545 ;
        RECT 109.290 201.125 109.550 201.445 ;
        RECT 108.815 200.950 109.115 201.015 ;
        RECT 108.805 200.690 109.125 200.950 ;
        RECT 108.815 200.625 109.115 200.690 ;
        RECT 108.815 189.145 109.115 189.210 ;
        RECT 108.805 188.885 109.125 189.145 ;
        RECT 108.815 188.820 109.115 188.885 ;
        RECT 108.805 186.430 109.125 186.475 ;
        RECT 109.335 186.430 109.505 201.125 ;
        RECT 108.805 186.260 109.505 186.430 ;
        RECT 108.805 186.215 109.125 186.260 ;
        RECT 109.790 185.965 109.960 201.545 ;
        RECT 110.790 201.125 111.050 201.445 ;
        RECT 110.315 200.950 110.615 201.015 ;
        RECT 110.305 200.690 110.625 200.950 ;
        RECT 110.315 200.625 110.615 200.690 ;
        RECT 110.315 189.145 110.615 189.210 ;
        RECT 110.305 188.885 110.625 189.145 ;
        RECT 110.315 188.820 110.615 188.885 ;
        RECT 110.305 186.430 110.625 186.475 ;
        RECT 110.835 186.430 111.005 201.125 ;
        RECT 110.305 186.260 111.005 186.430 ;
        RECT 110.305 186.215 110.625 186.260 ;
        RECT 111.290 185.965 111.460 201.545 ;
        RECT 112.290 201.125 112.550 201.445 ;
        RECT 111.815 200.950 112.115 201.015 ;
        RECT 111.805 200.690 112.125 200.950 ;
        RECT 111.815 200.625 112.115 200.690 ;
        RECT 111.815 189.145 112.115 189.210 ;
        RECT 111.805 188.885 112.125 189.145 ;
        RECT 111.815 188.820 112.115 188.885 ;
        RECT 111.805 186.430 112.125 186.475 ;
        RECT 112.335 186.430 112.505 201.125 ;
        RECT 111.805 186.260 112.505 186.430 ;
        RECT 111.805 186.215 112.125 186.260 ;
        RECT 112.790 185.965 112.960 201.545 ;
        RECT 113.790 201.125 114.050 201.445 ;
        RECT 113.315 200.950 113.615 201.015 ;
        RECT 113.305 200.690 113.625 200.950 ;
        RECT 113.315 200.625 113.615 200.690 ;
        RECT 113.315 189.145 113.615 189.210 ;
        RECT 113.305 188.885 113.625 189.145 ;
        RECT 113.315 188.820 113.615 188.885 ;
        RECT 113.305 186.430 113.625 186.475 ;
        RECT 113.835 186.430 114.005 201.125 ;
        RECT 113.305 186.260 114.005 186.430 ;
        RECT 113.305 186.215 113.625 186.260 ;
        RECT 114.290 185.965 114.460 201.545 ;
        RECT 115.290 201.125 115.550 201.445 ;
        RECT 114.815 200.950 115.115 201.015 ;
        RECT 114.805 200.690 115.125 200.950 ;
        RECT 114.815 200.625 115.115 200.690 ;
        RECT 114.815 189.145 115.115 189.210 ;
        RECT 114.805 188.885 115.125 189.145 ;
        RECT 114.815 188.820 115.115 188.885 ;
        RECT 114.805 186.430 115.125 186.475 ;
        RECT 115.335 186.430 115.505 201.125 ;
        RECT 114.805 186.260 115.505 186.430 ;
        RECT 114.805 186.215 115.125 186.260 ;
        RECT 115.790 185.965 115.960 201.545 ;
        RECT 116.790 201.125 117.050 201.445 ;
        RECT 116.315 200.950 116.615 201.015 ;
        RECT 116.305 200.690 116.625 200.950 ;
        RECT 116.315 200.625 116.615 200.690 ;
        RECT 116.315 189.145 116.615 189.210 ;
        RECT 116.305 188.885 116.625 189.145 ;
        RECT 116.315 188.820 116.615 188.885 ;
        RECT 116.305 186.430 116.625 186.475 ;
        RECT 116.835 186.430 117.005 201.125 ;
        RECT 116.305 186.260 117.005 186.430 ;
        RECT 116.305 186.215 116.625 186.260 ;
        RECT 117.290 185.965 117.460 201.545 ;
        RECT 118.290 201.125 118.550 201.445 ;
        RECT 117.815 200.950 118.115 201.015 ;
        RECT 117.805 200.690 118.125 200.950 ;
        RECT 117.815 200.625 118.115 200.690 ;
        RECT 117.815 189.145 118.115 189.210 ;
        RECT 117.805 188.885 118.125 189.145 ;
        RECT 117.815 188.820 118.115 188.885 ;
        RECT 117.805 186.430 118.125 186.475 ;
        RECT 118.335 186.430 118.505 201.125 ;
        RECT 117.805 186.260 118.505 186.430 ;
        RECT 117.805 186.215 118.125 186.260 ;
        RECT 118.790 185.965 118.960 201.545 ;
        RECT 119.435 200.965 119.735 201.015 ;
        RECT 119.410 200.675 119.760 200.965 ;
        RECT 119.435 200.625 119.735 200.675 ;
        RECT 119.285 189.160 119.585 189.210 ;
        RECT 119.260 188.870 119.610 189.160 ;
        RECT 119.285 188.820 119.585 188.870 ;
        RECT 107.380 185.795 108.460 185.965 ;
        RECT 108.880 185.795 109.960 185.965 ;
        RECT 110.380 185.795 111.460 185.965 ;
        RECT 111.880 185.795 112.960 185.965 ;
        RECT 113.380 185.795 114.460 185.965 ;
        RECT 114.880 185.795 115.960 185.965 ;
        RECT 116.380 185.795 117.460 185.965 ;
        RECT 117.880 185.795 118.960 185.965 ;
        RECT 76.725 183.940 77.025 184.005 ;
        RECT 76.715 183.680 77.035 183.940 ;
        RECT 76.725 183.615 77.025 183.680 ;
        RECT 77.385 183.615 77.685 184.005 ;
        RECT 106.630 183.530 106.980 183.575 ;
        RECT 76.290 183.185 76.550 183.505 ;
        RECT 106.600 183.180 107.010 183.530 ;
        RECT 106.630 183.135 106.980 183.180 ;
        RECT 39.335 182.765 39.595 183.085 ;
        RECT 40.835 182.765 41.095 183.085 ;
        RECT 42.335 182.765 42.595 183.085 ;
        RECT 43.835 182.765 44.095 183.085 ;
        RECT 45.335 182.765 45.595 183.085 ;
        RECT 46.835 182.765 47.095 183.085 ;
        RECT 48.335 182.765 48.595 183.085 ;
        RECT 49.835 182.765 50.095 183.085 ;
        RECT 65.335 182.765 65.595 183.085 ;
        RECT 66.835 182.765 67.095 183.085 ;
        RECT 68.335 182.765 68.595 183.085 ;
        RECT 69.835 182.765 70.095 183.085 ;
        RECT 71.335 182.765 71.595 183.085 ;
        RECT 72.835 182.765 73.095 183.085 ;
        RECT 74.335 182.765 74.595 183.085 ;
        RECT 75.835 182.765 76.095 183.085 ;
        RECT 106.730 182.480 107.080 182.525 ;
        RECT 106.700 182.130 107.110 182.480 ;
        RECT 106.730 182.085 107.080 182.130 ;
        RECT 107.380 179.295 107.550 185.795 ;
        RECT 107.790 185.265 108.050 185.585 ;
        RECT 107.835 181.485 108.005 185.265 ;
        RECT 108.215 184.110 108.535 184.370 ;
        RECT 108.290 182.045 108.460 184.110 ;
        RECT 108.290 181.800 108.600 182.045 ;
        RECT 108.340 181.725 108.600 181.800 ;
        RECT 108.245 181.485 108.505 181.560 ;
        RECT 107.835 181.315 108.505 181.485 ;
        RECT 108.245 181.240 108.505 181.315 ;
        RECT 108.880 179.295 109.050 185.795 ;
        RECT 109.290 185.265 109.550 185.585 ;
        RECT 109.335 181.485 109.505 185.265 ;
        RECT 109.715 184.110 110.035 184.370 ;
        RECT 109.790 182.045 109.960 184.110 ;
        RECT 109.790 181.800 110.100 182.045 ;
        RECT 109.840 181.725 110.100 181.800 ;
        RECT 109.745 181.485 110.005 181.560 ;
        RECT 109.335 181.315 110.005 181.485 ;
        RECT 109.745 181.240 110.005 181.315 ;
        RECT 110.380 179.295 110.550 185.795 ;
        RECT 110.790 185.265 111.050 185.585 ;
        RECT 110.835 181.485 111.005 185.265 ;
        RECT 111.215 184.110 111.535 184.370 ;
        RECT 111.290 182.045 111.460 184.110 ;
        RECT 111.290 181.800 111.600 182.045 ;
        RECT 111.340 181.725 111.600 181.800 ;
        RECT 111.245 181.485 111.505 181.560 ;
        RECT 110.835 181.315 111.505 181.485 ;
        RECT 111.245 181.240 111.505 181.315 ;
        RECT 111.880 179.295 112.050 185.795 ;
        RECT 112.290 185.265 112.550 185.585 ;
        RECT 112.335 181.485 112.505 185.265 ;
        RECT 112.715 184.110 113.035 184.370 ;
        RECT 112.790 182.045 112.960 184.110 ;
        RECT 112.790 181.800 113.100 182.045 ;
        RECT 112.840 181.725 113.100 181.800 ;
        RECT 112.745 181.485 113.005 181.560 ;
        RECT 112.335 181.315 113.005 181.485 ;
        RECT 112.745 181.240 113.005 181.315 ;
        RECT 113.380 179.295 113.550 185.795 ;
        RECT 113.790 185.265 114.050 185.585 ;
        RECT 113.835 181.485 114.005 185.265 ;
        RECT 114.215 184.110 114.535 184.370 ;
        RECT 114.290 182.045 114.460 184.110 ;
        RECT 114.290 181.800 114.600 182.045 ;
        RECT 114.340 181.725 114.600 181.800 ;
        RECT 114.245 181.485 114.505 181.560 ;
        RECT 113.835 181.315 114.505 181.485 ;
        RECT 114.245 181.240 114.505 181.315 ;
        RECT 114.880 179.295 115.050 185.795 ;
        RECT 115.290 185.265 115.550 185.585 ;
        RECT 115.335 181.485 115.505 185.265 ;
        RECT 115.715 184.110 116.035 184.370 ;
        RECT 115.790 182.045 115.960 184.110 ;
        RECT 115.790 181.800 116.100 182.045 ;
        RECT 115.840 181.725 116.100 181.800 ;
        RECT 115.745 181.485 116.005 181.560 ;
        RECT 115.335 181.315 116.005 181.485 ;
        RECT 115.745 181.240 116.005 181.315 ;
        RECT 116.380 179.295 116.550 185.795 ;
        RECT 116.790 185.265 117.050 185.585 ;
        RECT 116.835 181.485 117.005 185.265 ;
        RECT 117.215 184.110 117.535 184.370 ;
        RECT 117.290 182.045 117.460 184.110 ;
        RECT 117.290 181.800 117.600 182.045 ;
        RECT 117.340 181.725 117.600 181.800 ;
        RECT 117.245 181.485 117.505 181.560 ;
        RECT 116.835 181.315 117.505 181.485 ;
        RECT 117.245 181.240 117.505 181.315 ;
        RECT 117.880 179.295 118.050 185.795 ;
        RECT 118.290 185.265 118.550 185.585 ;
        RECT 118.335 181.485 118.505 185.265 ;
        RECT 118.715 184.110 119.035 184.370 ;
        RECT 118.790 182.045 118.960 184.110 ;
        RECT 119.410 183.530 119.760 183.575 ;
        RECT 119.380 183.180 119.790 183.530 ;
        RECT 119.410 183.135 119.760 183.180 ;
        RECT 119.265 182.480 119.615 182.525 ;
        RECT 119.235 182.130 119.645 182.480 ;
        RECT 119.265 182.085 119.615 182.130 ;
        RECT 118.790 181.800 119.100 182.045 ;
        RECT 118.840 181.725 119.100 181.800 ;
        RECT 118.745 181.485 119.005 181.560 ;
        RECT 118.335 181.315 119.005 181.485 ;
        RECT 118.745 181.240 119.005 181.315 ;
        RECT 107.380 179.125 108.005 179.295 ;
        RECT 108.880 179.125 109.505 179.295 ;
        RECT 110.380 179.125 111.005 179.295 ;
        RECT 111.880 179.125 112.505 179.295 ;
        RECT 113.380 179.125 114.005 179.295 ;
        RECT 114.880 179.125 115.505 179.295 ;
        RECT 116.380 179.125 117.005 179.295 ;
        RECT 117.880 179.125 118.505 179.295 ;
        RECT 38.755 178.295 39.055 178.345 ;
        RECT 38.730 178.005 39.080 178.295 ;
        RECT 38.755 177.955 39.055 178.005 ;
        RECT 39.745 171.845 40.095 178.830 ;
        RECT 40.295 178.280 40.595 178.345 ;
        RECT 40.285 178.020 40.605 178.280 ;
        RECT 40.295 177.955 40.595 178.020 ;
        RECT 38.595 171.495 40.095 171.845 ;
        RECT 38.595 167.845 38.945 171.495 ;
        RECT 41.245 170.845 41.595 178.830 ;
        RECT 41.795 178.280 42.095 178.345 ;
        RECT 41.785 178.020 42.105 178.280 ;
        RECT 41.795 177.955 42.095 178.020 ;
        RECT 40.875 170.495 41.595 170.845 ;
        RECT 38.565 167.495 38.975 167.845 ;
        RECT 40.875 166.845 41.225 170.495 ;
        RECT 42.745 169.845 43.095 178.830 ;
        RECT 43.295 178.280 43.595 178.345 ;
        RECT 43.285 178.020 43.605 178.280 ;
        RECT 43.295 177.955 43.595 178.020 ;
        RECT 44.245 169.845 44.595 178.830 ;
        RECT 44.795 178.280 45.095 178.345 ;
        RECT 44.785 178.020 45.105 178.280 ;
        RECT 44.795 177.955 45.095 178.020 ;
        RECT 45.745 169.845 46.095 178.830 ;
        RECT 46.295 178.280 46.595 178.345 ;
        RECT 46.285 178.020 46.605 178.280 ;
        RECT 46.295 177.955 46.595 178.020 ;
        RECT 41.950 169.495 43.095 169.845 ;
        RECT 44.230 169.495 44.595 169.845 ;
        RECT 45.305 169.495 46.095 169.845 ;
        RECT 47.245 169.845 47.595 178.830 ;
        RECT 47.795 178.280 48.095 178.345 ;
        RECT 47.785 178.020 48.105 178.280 ;
        RECT 47.795 177.955 48.095 178.020 ;
        RECT 48.745 169.845 49.095 178.830 ;
        RECT 49.295 178.280 49.595 178.345 ;
        RECT 49.285 178.020 49.605 178.280 ;
        RECT 49.295 177.955 49.595 178.020 ;
        RECT 47.245 169.495 47.935 169.845 ;
        RECT 40.845 166.495 41.255 166.845 ;
        RECT 41.950 165.845 42.300 169.495 ;
        RECT 43.125 167.495 43.535 167.845 ;
        RECT 39.640 165.495 40.050 165.845 ;
        RECT 41.920 165.495 42.330 165.845 ;
        RECT 29.705 159.495 30.115 159.845 ;
        RECT 26.220 157.495 26.630 157.845 ;
        RECT 26.250 148.135 26.600 157.495 ;
        RECT 29.735 148.135 30.085 159.495 ;
        RECT 36.415 155.495 36.825 155.845 ;
        RECT 32.930 153.495 33.340 153.845 ;
        RECT 32.960 148.135 33.310 153.495 ;
        RECT 36.445 148.135 36.795 155.495 ;
        RECT 39.670 148.135 40.020 165.495 ;
        RECT 43.155 148.135 43.505 167.495 ;
        RECT 44.230 164.845 44.580 169.495 ;
        RECT 44.200 164.495 44.610 164.845 ;
        RECT 45.305 163.845 45.655 169.495 ;
        RECT 45.275 163.495 45.685 163.845 ;
        RECT 47.585 162.845 47.935 169.495 ;
        RECT 48.660 169.495 49.095 169.845 ;
        RECT 50.245 169.845 50.595 178.830 ;
        RECT 50.795 178.280 51.095 178.345 ;
        RECT 51.285 178.295 51.585 178.345 ;
        RECT 64.755 178.295 65.055 178.345 ;
        RECT 50.785 178.020 51.105 178.280 ;
        RECT 50.795 177.955 51.095 178.020 ;
        RECT 51.260 178.005 51.610 178.295 ;
        RECT 64.730 178.005 65.080 178.295 ;
        RECT 51.285 177.955 51.585 178.005 ;
        RECT 64.755 177.955 65.055 178.005 ;
        RECT 65.745 169.845 66.095 178.830 ;
        RECT 66.295 178.280 66.595 178.345 ;
        RECT 66.285 178.020 66.605 178.280 ;
        RECT 66.295 177.955 66.595 178.020 ;
        RECT 50.245 169.495 51.290 169.845 ;
        RECT 47.555 162.495 47.965 162.845 ;
        RECT 48.660 161.845 49.010 169.495 ;
        RECT 49.835 163.495 50.245 163.845 ;
        RECT 46.350 161.495 46.760 161.845 ;
        RECT 48.630 161.495 49.040 161.845 ;
        RECT 46.380 148.135 46.730 161.495 ;
        RECT 49.865 148.135 50.215 163.495 ;
        RECT 50.940 160.845 51.290 169.495 ;
        RECT 65.435 169.495 66.095 169.845 ;
        RECT 67.245 169.845 67.595 178.830 ;
        RECT 67.795 178.280 68.095 178.345 ;
        RECT 67.785 178.020 68.105 178.280 ;
        RECT 67.795 177.955 68.095 178.020 ;
        RECT 68.745 169.845 69.095 178.830 ;
        RECT 69.295 178.280 69.595 178.345 ;
        RECT 69.285 178.020 69.605 178.280 ;
        RECT 69.295 177.955 69.595 178.020 ;
        RECT 70.245 169.845 70.595 178.830 ;
        RECT 70.795 178.280 71.095 178.345 ;
        RECT 70.785 178.020 71.105 178.280 ;
        RECT 70.795 177.955 71.095 178.020 ;
        RECT 71.745 170.845 72.095 178.830 ;
        RECT 72.295 178.280 72.595 178.345 ;
        RECT 72.285 178.020 72.605 178.280 ;
        RECT 72.295 177.955 72.595 178.020 ;
        RECT 71.745 170.495 72.495 170.845 ;
        RECT 67.245 169.495 68.065 169.845 ;
        RECT 68.745 169.495 69.140 169.845 ;
        RECT 70.245 169.495 71.420 169.845 ;
        RECT 50.910 160.495 51.320 160.845 ;
        RECT 65.435 159.845 65.785 169.495 ;
        RECT 66.480 164.495 66.890 164.845 ;
        RECT 65.405 159.495 65.815 159.845 ;
        RECT 56.545 158.495 56.955 158.845 ;
        RECT 53.060 156.495 53.470 156.845 ;
        RECT 53.090 148.135 53.440 156.495 ;
        RECT 56.575 148.135 56.925 158.495 ;
        RECT 63.255 154.495 63.665 154.845 ;
        RECT 59.770 152.495 60.180 152.845 ;
        RECT 59.800 148.135 60.150 152.495 ;
        RECT 63.285 148.135 63.635 154.495 ;
        RECT 66.510 148.135 66.860 164.495 ;
        RECT 67.715 158.845 68.065 169.495 ;
        RECT 67.685 158.495 68.095 158.845 ;
        RECT 68.790 157.845 69.140 169.495 ;
        RECT 69.965 166.495 70.375 166.845 ;
        RECT 68.760 157.495 69.170 157.845 ;
        RECT 69.995 148.135 70.345 166.495 ;
        RECT 71.070 156.845 71.420 169.495 ;
        RECT 71.040 156.495 71.450 156.845 ;
        RECT 72.145 155.845 72.495 170.495 ;
        RECT 73.245 169.845 73.595 178.830 ;
        RECT 73.795 178.280 74.095 178.345 ;
        RECT 73.785 178.020 74.105 178.280 ;
        RECT 73.795 177.955 74.095 178.020 ;
        RECT 74.745 170.845 75.095 178.830 ;
        RECT 75.295 178.280 75.595 178.345 ;
        RECT 75.285 178.020 75.605 178.280 ;
        RECT 75.295 177.955 75.595 178.020 ;
        RECT 76.245 171.845 76.595 178.830 ;
        RECT 107.835 178.440 108.005 179.125 ;
        RECT 109.335 178.440 109.505 179.125 ;
        RECT 110.835 178.440 111.005 179.125 ;
        RECT 112.335 178.440 112.505 179.125 ;
        RECT 113.835 178.440 114.005 179.125 ;
        RECT 115.335 178.440 115.505 179.125 ;
        RECT 116.835 178.440 117.005 179.125 ;
        RECT 118.335 178.440 118.505 179.125 ;
        RECT 76.795 178.280 77.095 178.345 ;
        RECT 77.285 178.295 77.585 178.345 ;
        RECT 76.785 178.020 77.105 178.280 ;
        RECT 76.795 177.955 77.095 178.020 ;
        RECT 77.260 178.005 77.610 178.295 ;
        RECT 107.760 178.180 108.080 178.440 ;
        RECT 109.260 178.180 109.580 178.440 ;
        RECT 110.760 178.180 111.080 178.440 ;
        RECT 112.260 178.180 112.580 178.440 ;
        RECT 113.760 178.180 114.080 178.440 ;
        RECT 115.260 178.180 115.580 178.440 ;
        RECT 116.760 178.180 117.080 178.440 ;
        RECT 118.260 178.180 118.580 178.440 ;
        RECT 77.285 177.955 77.585 178.005 ;
        RECT 106.655 176.790 106.955 176.840 ;
        RECT 106.630 176.500 106.980 176.790 ;
        RECT 107.310 176.775 107.610 176.840 ;
        RECT 107.300 176.515 107.620 176.775 ;
        RECT 106.655 176.450 106.955 176.500 ;
        RECT 107.310 176.450 107.610 176.515 ;
        RECT 76.245 171.495 78.130 171.845 ;
        RECT 74.745 170.495 75.850 170.845 ;
        RECT 73.245 169.495 74.775 169.845 ;
        RECT 73.190 160.495 73.600 160.845 ;
        RECT 72.115 155.495 72.525 155.845 ;
        RECT 73.220 148.135 73.570 160.495 ;
        RECT 74.425 154.845 74.775 169.495 ;
        RECT 74.395 154.495 74.805 154.845 ;
        RECT 75.500 153.845 75.850 170.495 ;
        RECT 76.675 162.495 77.085 162.845 ;
        RECT 75.470 153.495 75.880 153.845 ;
        RECT 76.705 148.135 77.055 162.495 ;
        RECT 77.780 152.845 78.130 171.495 ;
        RECT 77.750 152.495 78.160 152.845 ;
        RECT 26.340 142.270 26.510 148.135 ;
        RECT 29.825 146.770 29.995 148.135 ;
        RECT 29.715 146.470 30.105 146.770 ;
        RECT 27.595 146.035 27.915 146.295 ;
        RECT 26.710 145.720 27.100 146.020 ;
        RECT 26.710 142.720 27.100 143.020 ;
        RECT 26.230 141.970 26.620 142.270 ;
        RECT 27.670 141.795 27.840 146.035 ;
        RECT 29.825 145.250 29.995 146.470 ;
        RECT 29.750 144.990 30.070 145.250 ;
        RECT 28.435 144.535 28.755 144.795 ;
        RECT 27.595 141.535 27.915 141.795 ;
        RECT 26.710 139.720 27.100 140.020 ;
        RECT 26.710 136.720 27.100 137.020 ;
        RECT 27.670 134.770 27.840 141.535 ;
        RECT 28.015 140.035 28.335 140.295 ;
        RECT 28.090 137.770 28.260 140.035 ;
        RECT 27.980 137.470 28.370 137.770 ;
        RECT 28.510 136.270 28.680 144.535 ;
        RECT 29.825 143.750 29.995 144.990 ;
        RECT 32.370 144.220 32.760 144.520 ;
        RECT 29.750 143.490 30.070 143.750 ;
        RECT 28.855 143.035 29.175 143.295 ;
        RECT 28.930 138.795 29.100 143.035 ;
        RECT 33.050 142.270 33.220 148.135 ;
        RECT 36.535 146.770 36.705 148.135 ;
        RECT 36.425 146.470 36.815 146.770 ;
        RECT 34.305 146.035 34.625 146.295 ;
        RECT 33.420 145.720 33.810 146.020 ;
        RECT 33.420 142.720 33.810 143.020 ;
        RECT 29.715 141.970 30.105 142.270 ;
        RECT 32.940 141.970 33.330 142.270 ;
        RECT 29.825 140.750 29.995 141.970 ;
        RECT 34.380 141.795 34.550 146.035 ;
        RECT 36.535 145.250 36.705 146.470 ;
        RECT 36.460 144.990 36.780 145.250 ;
        RECT 35.145 144.535 35.465 144.795 ;
        RECT 34.305 141.535 34.625 141.795 ;
        RECT 32.370 141.220 32.760 141.520 ;
        RECT 29.750 140.490 30.070 140.750 ;
        RECT 29.825 139.250 29.995 140.490 ;
        RECT 33.420 139.720 33.810 140.020 ;
        RECT 29.750 138.990 30.070 139.250 ;
        RECT 31.520 138.970 31.910 139.270 ;
        RECT 28.855 138.535 29.175 138.795 ;
        RECT 28.930 136.655 29.100 138.535 ;
        RECT 31.630 137.750 31.800 138.970 ;
        RECT 32.370 138.220 32.760 138.520 ;
        RECT 31.555 137.490 31.875 137.750 ;
        RECT 29.750 137.035 30.070 137.295 ;
        RECT 28.860 136.395 29.180 136.655 ;
        RECT 28.400 135.970 28.790 136.270 ;
        RECT 28.930 136.035 29.100 136.395 ;
        RECT 29.825 136.250 29.995 137.035 ;
        RECT 33.420 136.720 33.810 137.020 ;
        RECT 29.750 135.990 30.070 136.250 ;
        RECT 29.780 135.505 30.040 135.825 ;
        RECT 27.560 134.470 27.950 134.770 ;
        RECT 26.710 133.720 27.100 134.020 ;
        RECT 29.825 132.135 29.995 135.505 ;
        RECT 32.370 135.220 32.760 135.520 ;
        RECT 34.380 134.770 34.550 141.535 ;
        RECT 34.725 140.035 35.045 140.295 ;
        RECT 34.800 137.770 34.970 140.035 ;
        RECT 34.690 137.470 35.080 137.770 ;
        RECT 35.220 136.270 35.390 144.535 ;
        RECT 36.535 143.750 36.705 144.990 ;
        RECT 39.080 144.220 39.470 144.520 ;
        RECT 36.460 143.490 36.780 143.750 ;
        RECT 35.565 143.035 35.885 143.295 ;
        RECT 35.640 139.315 35.810 143.035 ;
        RECT 39.760 142.270 39.930 148.135 ;
        RECT 43.245 146.770 43.415 148.135 ;
        RECT 43.135 146.470 43.525 146.770 ;
        RECT 41.015 146.035 41.335 146.295 ;
        RECT 40.130 145.720 40.520 146.020 ;
        RECT 40.130 142.720 40.520 143.020 ;
        RECT 36.425 141.970 36.815 142.270 ;
        RECT 39.650 141.970 40.040 142.270 ;
        RECT 36.535 140.750 36.705 141.970 ;
        RECT 41.090 141.795 41.260 146.035 ;
        RECT 43.245 145.250 43.415 146.470 ;
        RECT 43.170 144.990 43.490 145.250 ;
        RECT 41.855 144.535 42.175 144.795 ;
        RECT 41.015 141.535 41.335 141.795 ;
        RECT 39.080 141.220 39.470 141.520 ;
        RECT 36.460 140.490 36.780 140.750 ;
        RECT 35.575 138.795 35.875 139.315 ;
        RECT 36.535 139.250 36.705 140.490 ;
        RECT 40.130 139.720 40.520 140.020 ;
        RECT 36.460 138.990 36.780 139.250 ;
        RECT 35.565 138.535 35.885 138.795 ;
        RECT 35.640 137.535 35.810 138.535 ;
        RECT 39.080 138.220 39.470 138.520 ;
        RECT 36.460 137.035 36.780 137.295 ;
        RECT 35.110 135.970 35.500 136.270 ;
        RECT 36.535 136.250 36.705 137.035 ;
        RECT 40.130 136.720 40.520 137.020 ;
        RECT 36.460 135.990 36.780 136.250 ;
        RECT 36.490 135.505 36.750 135.825 ;
        RECT 34.270 134.470 34.660 134.770 ;
        RECT 33.420 133.720 33.810 134.020 ;
        RECT 29.750 131.875 30.070 132.135 ;
        RECT 36.535 131.750 36.705 135.505 ;
        RECT 39.080 135.220 39.470 135.520 ;
        RECT 41.090 134.770 41.260 141.535 ;
        RECT 41.435 140.035 41.755 140.295 ;
        RECT 41.510 137.770 41.680 140.035 ;
        RECT 41.400 137.470 41.790 137.770 ;
        RECT 41.930 136.270 42.100 144.535 ;
        RECT 43.245 143.750 43.415 144.990 ;
        RECT 45.790 144.220 46.180 144.520 ;
        RECT 43.170 143.490 43.490 143.750 ;
        RECT 42.275 143.035 42.595 143.295 ;
        RECT 42.350 138.795 42.520 143.035 ;
        RECT 46.470 142.270 46.640 148.135 ;
        RECT 49.955 146.770 50.125 148.135 ;
        RECT 49.845 146.470 50.235 146.770 ;
        RECT 47.725 146.035 48.045 146.295 ;
        RECT 46.840 145.720 47.230 146.020 ;
        RECT 46.840 142.720 47.230 143.020 ;
        RECT 43.135 141.970 43.525 142.270 ;
        RECT 46.360 141.970 46.750 142.270 ;
        RECT 43.245 140.750 43.415 141.970 ;
        RECT 47.800 141.795 47.970 146.035 ;
        RECT 49.955 145.250 50.125 146.470 ;
        RECT 49.880 144.990 50.200 145.250 ;
        RECT 48.565 144.535 48.885 144.795 ;
        RECT 47.725 141.535 48.045 141.795 ;
        RECT 45.790 141.220 46.180 141.520 ;
        RECT 43.170 140.490 43.490 140.750 ;
        RECT 43.245 139.250 43.415 140.490 ;
        RECT 46.840 139.720 47.230 140.020 ;
        RECT 43.170 138.990 43.490 139.250 ;
        RECT 44.940 138.970 45.330 139.270 ;
        RECT 42.275 138.535 42.595 138.795 ;
        RECT 42.350 136.655 42.520 138.535 ;
        RECT 45.050 137.750 45.220 138.970 ;
        RECT 45.790 138.220 46.180 138.520 ;
        RECT 44.975 137.490 45.295 137.750 ;
        RECT 43.170 137.035 43.490 137.295 ;
        RECT 42.280 136.395 42.600 136.655 ;
        RECT 41.820 135.970 42.210 136.270 ;
        RECT 42.350 136.035 42.520 136.395 ;
        RECT 43.245 136.250 43.415 137.035 ;
        RECT 46.840 136.720 47.230 137.020 ;
        RECT 43.170 135.990 43.490 136.250 ;
        RECT 43.200 135.505 43.460 135.825 ;
        RECT 40.980 134.470 41.370 134.770 ;
        RECT 38.265 134.035 38.585 134.295 ;
        RECT 38.340 133.290 38.510 134.035 ;
        RECT 40.130 133.720 40.520 134.020 ;
        RECT 38.265 133.030 38.585 133.290 ;
        RECT 43.245 132.135 43.415 135.505 ;
        RECT 45.790 135.220 46.180 135.520 ;
        RECT 47.800 134.770 47.970 141.535 ;
        RECT 48.145 140.035 48.465 140.295 ;
        RECT 48.220 137.770 48.390 140.035 ;
        RECT 48.110 137.470 48.500 137.770 ;
        RECT 48.640 136.270 48.810 144.535 ;
        RECT 49.955 143.750 50.125 144.990 ;
        RECT 52.500 144.220 52.890 144.520 ;
        RECT 49.880 143.490 50.200 143.750 ;
        RECT 48.985 143.035 49.305 143.295 ;
        RECT 49.060 139.315 49.230 143.035 ;
        RECT 53.180 142.270 53.350 148.135 ;
        RECT 56.665 146.770 56.835 148.135 ;
        RECT 56.555 146.470 56.945 146.770 ;
        RECT 54.435 146.035 54.755 146.295 ;
        RECT 53.550 145.720 53.940 146.020 ;
        RECT 53.550 142.720 53.940 143.020 ;
        RECT 49.845 141.970 50.235 142.270 ;
        RECT 53.070 141.970 53.460 142.270 ;
        RECT 49.955 140.750 50.125 141.970 ;
        RECT 54.510 141.795 54.680 146.035 ;
        RECT 56.665 145.250 56.835 146.470 ;
        RECT 56.590 144.990 56.910 145.250 ;
        RECT 55.275 144.535 55.595 144.795 ;
        RECT 54.435 141.535 54.755 141.795 ;
        RECT 52.500 141.220 52.890 141.520 ;
        RECT 49.880 140.490 50.200 140.750 ;
        RECT 48.995 138.795 49.295 139.315 ;
        RECT 49.955 139.250 50.125 140.490 ;
        RECT 53.550 139.720 53.940 140.020 ;
        RECT 49.880 138.990 50.200 139.250 ;
        RECT 48.985 138.535 49.305 138.795 ;
        RECT 49.060 137.535 49.230 138.535 ;
        RECT 52.500 138.220 52.890 138.520 ;
        RECT 49.880 137.035 50.200 137.295 ;
        RECT 48.530 135.970 48.920 136.270 ;
        RECT 49.955 136.250 50.125 137.035 ;
        RECT 53.550 136.720 53.940 137.020 ;
        RECT 49.880 135.990 50.200 136.250 ;
        RECT 49.910 135.505 50.170 135.825 ;
        RECT 47.690 134.470 48.080 134.770 ;
        RECT 46.840 133.720 47.230 134.020 ;
        RECT 43.170 131.875 43.490 132.135 ;
        RECT 49.955 131.750 50.125 135.505 ;
        RECT 52.500 135.220 52.890 135.520 ;
        RECT 54.510 134.770 54.680 141.535 ;
        RECT 54.855 140.035 55.175 140.295 ;
        RECT 54.930 137.770 55.100 140.035 ;
        RECT 54.820 137.470 55.210 137.770 ;
        RECT 55.350 136.270 55.520 144.535 ;
        RECT 56.665 143.750 56.835 144.990 ;
        RECT 59.210 144.220 59.600 144.520 ;
        RECT 56.590 143.490 56.910 143.750 ;
        RECT 55.695 143.035 56.015 143.295 ;
        RECT 55.770 138.795 55.940 143.035 ;
        RECT 59.890 142.270 60.060 148.135 ;
        RECT 63.375 146.770 63.545 148.135 ;
        RECT 63.265 146.470 63.655 146.770 ;
        RECT 61.145 146.035 61.465 146.295 ;
        RECT 60.260 145.720 60.650 146.020 ;
        RECT 60.260 142.720 60.650 143.020 ;
        RECT 56.555 141.970 56.945 142.270 ;
        RECT 59.780 141.970 60.170 142.270 ;
        RECT 56.665 140.750 56.835 141.970 ;
        RECT 61.220 141.795 61.390 146.035 ;
        RECT 63.375 145.250 63.545 146.470 ;
        RECT 63.300 144.990 63.620 145.250 ;
        RECT 61.985 144.535 62.305 144.795 ;
        RECT 61.145 141.535 61.465 141.795 ;
        RECT 59.210 141.220 59.600 141.520 ;
        RECT 56.590 140.490 56.910 140.750 ;
        RECT 56.665 139.250 56.835 140.490 ;
        RECT 60.260 139.720 60.650 140.020 ;
        RECT 56.590 138.990 56.910 139.250 ;
        RECT 58.360 138.970 58.750 139.270 ;
        RECT 55.695 138.535 56.015 138.795 ;
        RECT 55.770 136.655 55.940 138.535 ;
        RECT 58.470 137.750 58.640 138.970 ;
        RECT 59.210 138.220 59.600 138.520 ;
        RECT 58.395 137.490 58.715 137.750 ;
        RECT 56.590 137.035 56.910 137.295 ;
        RECT 55.700 136.395 56.020 136.655 ;
        RECT 55.240 135.970 55.630 136.270 ;
        RECT 55.770 136.035 55.940 136.395 ;
        RECT 56.665 136.250 56.835 137.035 ;
        RECT 60.260 136.720 60.650 137.020 ;
        RECT 56.590 135.990 56.910 136.250 ;
        RECT 56.620 135.505 56.880 135.825 ;
        RECT 54.400 134.470 54.790 134.770 ;
        RECT 51.685 134.035 52.005 134.295 ;
        RECT 51.760 132.905 51.930 134.035 ;
        RECT 53.550 133.720 53.940 134.020 ;
        RECT 51.685 132.645 52.005 132.905 ;
        RECT 56.665 132.165 56.835 135.505 ;
        RECT 59.210 135.220 59.600 135.520 ;
        RECT 61.220 134.770 61.390 141.535 ;
        RECT 61.565 140.035 61.885 140.295 ;
        RECT 61.640 137.770 61.810 140.035 ;
        RECT 61.530 137.470 61.920 137.770 ;
        RECT 62.060 136.270 62.230 144.535 ;
        RECT 63.375 143.750 63.545 144.990 ;
        RECT 65.920 144.220 66.310 144.520 ;
        RECT 63.300 143.490 63.620 143.750 ;
        RECT 62.405 143.035 62.725 143.295 ;
        RECT 62.480 139.315 62.650 143.035 ;
        RECT 66.600 142.270 66.770 148.135 ;
        RECT 70.085 146.770 70.255 148.135 ;
        RECT 69.975 146.470 70.365 146.770 ;
        RECT 67.855 146.035 68.175 146.295 ;
        RECT 66.970 145.720 67.360 146.020 ;
        RECT 66.970 142.720 67.360 143.020 ;
        RECT 63.265 141.970 63.655 142.270 ;
        RECT 66.490 141.970 66.880 142.270 ;
        RECT 63.375 140.750 63.545 141.970 ;
        RECT 67.930 141.795 68.100 146.035 ;
        RECT 70.085 145.250 70.255 146.470 ;
        RECT 70.010 144.990 70.330 145.250 ;
        RECT 68.695 144.535 69.015 144.795 ;
        RECT 67.855 141.535 68.175 141.795 ;
        RECT 65.920 141.220 66.310 141.520 ;
        RECT 63.300 140.490 63.620 140.750 ;
        RECT 62.415 138.795 62.715 139.315 ;
        RECT 63.375 139.250 63.545 140.490 ;
        RECT 66.970 139.720 67.360 140.020 ;
        RECT 63.300 138.990 63.620 139.250 ;
        RECT 62.405 138.535 62.725 138.795 ;
        RECT 62.480 137.535 62.650 138.535 ;
        RECT 65.920 138.220 66.310 138.520 ;
        RECT 63.300 137.035 63.620 137.295 ;
        RECT 61.950 135.970 62.340 136.270 ;
        RECT 63.375 136.250 63.545 137.035 ;
        RECT 66.970 136.720 67.360 137.020 ;
        RECT 63.300 135.990 63.620 136.250 ;
        RECT 63.330 135.505 63.590 135.825 ;
        RECT 61.110 134.470 61.500 134.770 ;
        RECT 60.260 133.720 60.650 134.020 ;
        RECT 56.620 131.845 56.880 132.165 ;
        RECT 63.375 131.750 63.545 135.505 ;
        RECT 65.920 135.220 66.310 135.520 ;
        RECT 67.930 134.770 68.100 141.535 ;
        RECT 68.275 140.035 68.595 140.295 ;
        RECT 68.350 137.770 68.520 140.035 ;
        RECT 68.240 137.470 68.630 137.770 ;
        RECT 68.770 136.270 68.940 144.535 ;
        RECT 70.085 143.750 70.255 144.990 ;
        RECT 72.630 144.220 73.020 144.520 ;
        RECT 70.010 143.490 70.330 143.750 ;
        RECT 69.115 143.035 69.435 143.295 ;
        RECT 69.190 138.795 69.360 143.035 ;
        RECT 73.310 142.270 73.480 148.135 ;
        RECT 76.795 146.770 76.965 148.135 ;
        RECT 76.685 146.470 77.075 146.770 ;
        RECT 83.395 146.470 83.785 146.770 ;
        RECT 90.105 146.470 90.495 146.770 ;
        RECT 74.565 146.035 74.885 146.295 ;
        RECT 73.680 145.720 74.070 146.020 ;
        RECT 73.680 142.720 74.070 143.020 ;
        RECT 69.975 141.970 70.365 142.270 ;
        RECT 73.200 141.970 73.590 142.270 ;
        RECT 70.085 140.750 70.255 141.970 ;
        RECT 74.640 141.795 74.810 146.035 ;
        RECT 76.795 145.250 76.965 146.470 ;
        RECT 81.275 146.035 81.595 146.295 ;
        RECT 80.390 145.720 80.780 146.020 ;
        RECT 76.720 144.990 77.040 145.250 ;
        RECT 75.405 144.535 75.725 144.795 ;
        RECT 74.565 141.535 74.885 141.795 ;
        RECT 72.630 141.220 73.020 141.520 ;
        RECT 70.010 140.490 70.330 140.750 ;
        RECT 70.085 139.250 70.255 140.490 ;
        RECT 73.680 139.720 74.070 140.020 ;
        RECT 70.010 138.990 70.330 139.250 ;
        RECT 71.780 138.970 72.170 139.270 ;
        RECT 69.115 138.535 69.435 138.795 ;
        RECT 69.190 136.655 69.360 138.535 ;
        RECT 71.890 137.750 72.060 138.970 ;
        RECT 72.630 138.220 73.020 138.520 ;
        RECT 71.815 137.490 72.135 137.750 ;
        RECT 70.010 137.035 70.330 137.295 ;
        RECT 69.120 136.395 69.440 136.655 ;
        RECT 68.660 135.970 69.050 136.270 ;
        RECT 69.190 136.035 69.360 136.395 ;
        RECT 70.085 136.250 70.255 137.035 ;
        RECT 73.680 136.720 74.070 137.020 ;
        RECT 70.010 135.990 70.330 136.250 ;
        RECT 70.040 135.505 70.300 135.825 ;
        RECT 67.820 134.470 68.210 134.770 ;
        RECT 65.105 134.035 65.425 134.295 ;
        RECT 65.180 132.520 65.350 134.035 ;
        RECT 66.970 133.720 67.360 134.020 ;
        RECT 65.105 132.260 65.425 132.520 ;
        RECT 70.085 132.135 70.255 135.505 ;
        RECT 72.630 135.220 73.020 135.520 ;
        RECT 74.640 134.770 74.810 141.535 ;
        RECT 74.985 140.035 75.305 140.295 ;
        RECT 75.060 137.770 75.230 140.035 ;
        RECT 74.950 137.470 75.340 137.770 ;
        RECT 75.480 136.270 75.650 144.535 ;
        RECT 76.795 143.750 76.965 144.990 ;
        RECT 79.340 144.220 79.730 144.520 ;
        RECT 76.720 143.490 77.040 143.750 ;
        RECT 75.825 143.035 76.145 143.295 ;
        RECT 75.900 139.315 76.070 143.035 ;
        RECT 80.390 142.720 80.780 143.020 ;
        RECT 76.685 141.970 77.075 142.270 ;
        RECT 79.910 141.970 80.300 142.270 ;
        RECT 76.795 140.750 76.965 141.970 ;
        RECT 79.340 141.220 79.730 141.520 ;
        RECT 76.720 140.490 77.040 140.750 ;
        RECT 75.835 138.795 76.135 139.315 ;
        RECT 76.795 139.250 76.965 140.490 ;
        RECT 76.720 138.990 77.040 139.250 ;
        RECT 75.825 138.535 76.145 138.795 ;
        RECT 75.900 137.535 76.070 138.535 ;
        RECT 79.340 138.220 79.730 138.520 ;
        RECT 76.720 137.035 77.040 137.295 ;
        RECT 75.370 135.970 75.760 136.270 ;
        RECT 76.795 136.250 76.965 137.035 ;
        RECT 76.720 135.990 77.040 136.250 ;
        RECT 76.750 135.505 77.010 135.825 ;
        RECT 74.530 134.470 74.920 134.770 ;
        RECT 73.680 133.720 74.070 134.020 ;
        RECT 70.010 131.875 70.330 132.135 ;
        RECT 36.460 131.490 36.780 131.750 ;
        RECT 49.880 131.490 50.200 131.750 ;
        RECT 63.300 131.490 63.620 131.750 ;
        RECT 70.085 131.420 70.255 131.875 ;
        RECT 76.795 131.750 76.965 135.505 ;
        RECT 79.340 135.220 79.730 135.520 ;
        RECT 78.525 134.035 78.845 134.295 ;
        RECT 78.600 132.135 78.770 134.035 ;
        RECT 80.020 132.905 80.190 141.970 ;
        RECT 81.350 141.795 81.520 146.035 ;
        RECT 83.505 145.250 83.675 146.470 ;
        RECT 87.985 146.035 88.305 146.295 ;
        RECT 87.100 145.720 87.490 146.020 ;
        RECT 83.430 144.990 83.750 145.250 ;
        RECT 82.115 144.535 82.435 144.795 ;
        RECT 81.275 141.535 81.595 141.795 ;
        RECT 80.390 139.720 80.780 140.020 ;
        RECT 80.390 136.720 80.780 137.020 ;
        RECT 81.350 134.770 81.520 141.535 ;
        RECT 81.695 140.035 82.015 140.295 ;
        RECT 81.770 137.770 81.940 140.035 ;
        RECT 81.660 137.470 82.050 137.770 ;
        RECT 82.190 136.270 82.360 144.535 ;
        RECT 83.505 143.750 83.675 144.990 ;
        RECT 86.050 144.220 86.440 144.520 ;
        RECT 83.430 143.705 83.750 143.750 ;
        RECT 83.085 143.535 83.750 143.705 ;
        RECT 82.535 143.035 82.855 143.295 ;
        RECT 82.610 138.795 82.780 143.035 ;
        RECT 82.535 138.535 82.855 138.795 ;
        RECT 82.610 136.655 82.780 138.535 ;
        RECT 82.540 136.395 82.860 136.655 ;
        RECT 82.080 135.970 82.470 136.270 ;
        RECT 82.610 136.035 82.780 136.395 ;
        RECT 81.240 134.470 81.630 134.770 ;
        RECT 80.390 133.720 80.780 134.020 ;
        RECT 83.085 133.290 83.255 143.535 ;
        RECT 83.430 143.490 83.750 143.535 ;
        RECT 87.100 142.720 87.490 143.020 ;
        RECT 83.395 141.970 83.785 142.270 ;
        RECT 86.620 141.970 87.010 142.270 ;
        RECT 83.505 140.750 83.675 141.970 ;
        RECT 86.050 141.220 86.440 141.520 ;
        RECT 83.430 140.490 83.750 140.750 ;
        RECT 83.505 139.250 83.675 140.490 ;
        RECT 83.430 138.990 83.750 139.250 ;
        RECT 85.200 138.970 85.590 139.270 ;
        RECT 85.310 137.750 85.480 138.970 ;
        RECT 86.050 138.220 86.440 138.520 ;
        RECT 85.235 137.490 85.555 137.750 ;
        RECT 83.430 137.035 83.750 137.295 ;
        RECT 83.505 136.250 83.675 137.035 ;
        RECT 83.430 135.990 83.750 136.250 ;
        RECT 83.460 135.505 83.720 135.825 ;
        RECT 83.010 133.030 83.330 133.290 ;
        RECT 79.945 132.645 80.265 132.905 ;
        RECT 78.525 131.875 78.845 132.135 ;
        RECT 76.720 131.490 77.040 131.750 ;
        RECT 69.995 123.645 70.345 131.420 ;
        RECT 69.965 123.295 70.375 123.645 ;
        RECT 76.705 122.145 77.055 131.490 ;
        RECT 83.505 131.410 83.675 135.505 ;
        RECT 86.050 135.220 86.440 135.520 ;
        RECT 86.730 132.135 86.900 141.970 ;
        RECT 88.060 141.795 88.230 146.035 ;
        RECT 90.215 145.250 90.385 146.470 ;
        RECT 90.140 144.990 90.460 145.250 ;
        RECT 88.825 144.535 89.145 144.795 ;
        RECT 87.985 141.535 88.305 141.795 ;
        RECT 87.100 139.720 87.490 140.020 ;
        RECT 87.100 136.720 87.490 137.020 ;
        RECT 88.060 134.770 88.230 141.535 ;
        RECT 88.405 140.035 88.725 140.295 ;
        RECT 88.480 137.770 88.650 140.035 ;
        RECT 88.370 137.470 88.760 137.770 ;
        RECT 88.900 136.270 89.070 144.535 ;
        RECT 90.215 143.750 90.385 144.990 ;
        RECT 92.760 144.220 93.150 144.520 ;
        RECT 90.140 143.705 90.460 143.750 ;
        RECT 89.795 143.535 90.460 143.705 ;
        RECT 89.245 143.035 89.565 143.295 ;
        RECT 89.320 139.315 89.490 143.035 ;
        RECT 89.255 138.795 89.555 139.315 ;
        RECT 89.245 138.535 89.565 138.795 ;
        RECT 89.320 137.535 89.490 138.535 ;
        RECT 88.790 135.970 89.180 136.270 ;
        RECT 87.950 134.470 88.340 134.770 ;
        RECT 87.100 133.720 87.490 134.020 ;
        RECT 89.795 132.520 89.965 143.535 ;
        RECT 90.140 143.490 90.460 143.535 ;
        RECT 90.105 141.970 90.495 142.270 ;
        RECT 90.215 140.750 90.385 141.970 ;
        RECT 92.760 141.220 93.150 141.520 ;
        RECT 90.140 140.490 90.460 140.750 ;
        RECT 90.215 139.250 90.385 140.490 ;
        RECT 90.140 138.990 90.460 139.250 ;
        RECT 92.760 138.220 93.150 138.520 ;
        RECT 90.140 137.035 90.460 137.295 ;
        RECT 90.215 136.250 90.385 137.035 ;
        RECT 90.140 135.990 90.460 136.250 ;
        RECT 90.170 135.505 90.430 135.825 ;
        RECT 89.720 132.260 90.040 132.520 ;
        RECT 86.655 131.875 86.975 132.135 ;
        RECT 90.215 131.435 90.385 135.505 ;
        RECT 92.760 135.220 93.150 135.520 ;
        RECT 91.945 134.035 92.265 134.295 ;
        RECT 92.020 133.290 92.190 134.035 ;
        RECT 91.945 133.030 92.265 133.290 ;
        RECT 76.675 121.795 77.085 122.145 ;
        RECT 83.415 120.645 83.765 131.410 ;
        RECT 90.125 125.145 90.475 131.435 ;
        RECT 90.095 124.795 90.505 125.145 ;
        RECT 108.200 124.750 108.550 177.705 ;
        RECT 108.810 176.775 109.110 176.840 ;
        RECT 108.800 176.515 109.120 176.775 ;
        RECT 108.810 176.450 109.110 176.515 ;
        RECT 109.700 123.250 110.050 177.705 ;
        RECT 110.310 176.775 110.610 176.840 ;
        RECT 110.300 176.515 110.620 176.775 ;
        RECT 110.310 176.450 110.610 176.515 ;
        RECT 111.200 121.750 111.550 177.705 ;
        RECT 111.810 176.775 112.110 176.840 ;
        RECT 111.800 176.515 112.120 176.775 ;
        RECT 111.810 176.450 112.110 176.515 ;
        RECT 74.320 120.295 74.730 120.645 ;
        RECT 83.385 120.295 83.795 120.645 ;
        RECT 15.980 118.795 16.390 119.145 ;
        RECT 16.010 37.445 16.360 118.795 ;
        RECT 17.480 117.295 17.890 117.645 ;
        RECT 17.510 57.575 17.860 117.295 ;
        RECT 18.980 115.795 19.390 116.145 ;
        RECT 17.480 57.225 17.890 57.575 ;
        RECT 19.010 50.865 19.360 115.795 ;
        RECT 20.480 114.295 20.890 114.645 ;
        RECT 18.980 50.515 19.390 50.865 ;
        RECT 20.510 44.155 20.860 114.295 ;
        RECT 42.025 101.230 42.325 101.340 ;
        RECT 42.025 101.060 47.320 101.230 ;
        RECT 42.025 100.950 42.325 101.060 ;
        RECT 33.775 100.470 34.075 100.860 ;
        RECT 36.775 100.470 37.075 100.860 ;
        RECT 39.775 100.470 40.075 100.860 ;
        RECT 42.775 100.470 43.075 100.860 ;
        RECT 45.775 100.470 46.075 100.860 ;
        RECT 34.525 99.900 34.825 100.010 ;
        RECT 41.590 99.900 41.850 99.975 ;
        RECT 46.090 99.900 46.350 99.975 ;
        RECT 34.525 99.730 46.350 99.900 ;
        RECT 34.525 99.620 34.825 99.730 ;
        RECT 41.590 99.655 41.850 99.730 ;
        RECT 46.090 99.655 46.350 99.730 ;
        RECT 37.525 99.480 37.825 99.590 ;
        RECT 40.090 99.480 40.350 99.555 ;
        RECT 37.525 99.310 40.350 99.480 ;
        RECT 37.525 99.200 37.825 99.310 ;
        RECT 40.090 99.235 40.350 99.310 ;
        RECT 36.025 99.060 36.325 99.170 ;
        RECT 44.590 99.060 44.850 99.135 ;
        RECT 36.025 98.890 44.850 99.060 ;
        RECT 36.025 98.780 36.325 98.890 ;
        RECT 44.590 98.815 44.850 98.890 ;
        RECT 36.450 98.640 36.710 98.710 ;
        RECT 38.590 98.640 38.850 98.715 ;
        RECT 43.090 98.640 43.350 98.715 ;
        RECT 36.090 98.470 43.350 98.640 ;
        RECT 36.450 98.390 36.710 98.470 ;
        RECT 38.590 98.395 38.850 98.470 ;
        RECT 43.090 98.395 43.350 98.470 ;
        RECT 47.150 98.375 47.320 101.060 ;
        RECT 47.150 98.205 48.020 98.375 ;
        RECT 31.930 97.745 32.190 97.820 ;
        RECT 35.560 97.745 35.880 97.790 ;
        RECT 31.930 97.575 35.880 97.745 ;
        RECT 31.930 97.500 32.190 97.575 ;
        RECT 35.560 97.530 35.880 97.575 ;
        RECT 36.045 97.745 36.305 97.820 ;
        RECT 37.090 97.745 37.350 97.820 ;
        RECT 36.045 97.575 37.350 97.745 ;
        RECT 36.045 97.500 36.305 97.575 ;
        RECT 37.090 97.500 37.350 97.575 ;
        RECT 39.045 97.745 39.305 97.820 ;
        RECT 40.545 97.745 40.805 97.820 ;
        RECT 42.025 97.745 42.325 97.855 ;
        RECT 39.045 97.575 42.325 97.745 ;
        RECT 39.045 97.500 39.305 97.575 ;
        RECT 40.545 97.500 40.805 97.575 ;
        RECT 42.025 97.465 42.325 97.575 ;
        RECT 43.545 97.745 43.805 97.820 ;
        RECT 45.045 97.745 45.305 97.820 ;
        RECT 46.525 97.745 46.825 97.855 ;
        RECT 43.545 97.575 47.390 97.745 ;
        RECT 43.545 97.500 43.805 97.575 ;
        RECT 45.045 97.500 45.305 97.575 ;
        RECT 46.525 97.465 46.825 97.575 ;
        RECT 47.220 96.420 47.390 97.575 ;
        RECT 47.850 97.050 48.020 98.205 ;
        RECT 48.415 97.050 48.715 97.160 ;
        RECT 47.850 96.880 48.715 97.050 ;
        RECT 48.415 96.770 48.715 96.880 ;
        RECT 49.045 96.420 49.345 96.530 ;
        RECT 47.220 96.250 49.345 96.420 ;
        RECT 49.045 96.140 49.345 96.250 ;
        RECT 65.655 96.060 66.345 99.915 ;
        RECT 37.545 95.940 37.805 96.015 ;
        RECT 39.025 95.940 39.325 96.050 ;
        RECT 37.545 95.770 39.325 95.940 ;
        RECT 37.545 95.695 37.805 95.770 ;
        RECT 39.025 95.660 39.325 95.770 ;
        RECT 54.480 95.370 69.155 96.060 ;
        RECT 35.275 94.810 35.575 95.200 ;
        RECT 38.275 94.810 38.575 95.200 ;
        RECT 41.275 94.810 41.575 95.200 ;
        RECT 44.275 94.810 44.575 95.200 ;
        RECT 42.025 94.520 42.325 94.630 ;
        RECT 47.155 94.520 47.455 94.630 ;
        RECT 42.025 94.350 47.455 94.520 ;
        RECT 54.480 94.500 55.170 95.370 ;
        RECT 42.025 94.240 42.325 94.350 ;
        RECT 47.155 94.240 47.455 94.350 ;
        RECT 33.775 93.760 34.075 94.150 ;
        RECT 36.775 93.760 37.075 94.150 ;
        RECT 39.775 93.760 40.075 94.150 ;
        RECT 42.775 93.760 43.075 94.150 ;
        RECT 45.775 93.760 46.075 94.150 ;
        RECT 54.450 93.810 55.200 94.500 ;
        RECT 56.045 94.285 56.735 94.975 ;
        RECT 57.425 94.285 58.115 94.975 ;
        RECT 58.805 94.285 59.495 94.975 ;
        RECT 60.185 94.285 60.875 94.975 ;
        RECT 61.565 94.285 62.255 94.975 ;
        RECT 62.945 94.285 63.635 94.975 ;
        RECT 64.325 94.285 65.015 94.975 ;
        RECT 65.705 94.285 66.395 94.975 ;
        RECT 67.085 94.285 67.775 94.975 ;
        RECT 68.465 94.285 69.155 94.975 ;
        RECT 55.535 93.725 56.365 94.045 ;
        RECT 34.525 93.190 34.825 93.300 ;
        RECT 41.590 93.190 41.850 93.265 ;
        RECT 46.090 93.190 46.350 93.265 ;
        RECT 34.525 93.020 46.350 93.190 ;
        RECT 34.525 92.910 34.825 93.020 ;
        RECT 41.590 92.945 41.850 93.020 ;
        RECT 46.090 92.945 46.350 93.020 ;
        RECT 55.535 93.070 56.250 93.725 ;
        RECT 56.505 93.530 56.735 94.285 ;
        RECT 56.915 93.725 57.745 94.045 ;
        RECT 56.505 93.210 56.765 93.530 ;
        RECT 56.915 93.355 57.630 93.725 ;
        RECT 57.400 93.070 57.630 93.355 ;
        RECT 57.885 93.530 58.115 94.285 ;
        RECT 58.295 93.725 59.125 94.045 ;
        RECT 57.885 93.210 58.145 93.530 ;
        RECT 58.295 93.355 59.010 93.725 ;
        RECT 58.780 93.070 59.010 93.355 ;
        RECT 59.265 93.530 59.495 94.285 ;
        RECT 59.675 93.725 60.505 94.045 ;
        RECT 59.265 93.210 59.525 93.530 ;
        RECT 59.675 93.355 60.390 93.725 ;
        RECT 60.160 93.070 60.390 93.355 ;
        RECT 60.645 93.530 60.875 94.285 ;
        RECT 61.055 93.725 61.885 94.045 ;
        RECT 60.645 93.210 60.905 93.530 ;
        RECT 61.055 93.355 61.770 93.725 ;
        RECT 61.540 93.070 61.770 93.355 ;
        RECT 62.025 93.530 62.255 94.285 ;
        RECT 62.435 93.725 63.265 94.045 ;
        RECT 62.025 93.210 62.285 93.530 ;
        RECT 62.435 93.355 63.150 93.725 ;
        RECT 62.920 93.070 63.150 93.355 ;
        RECT 63.405 93.530 63.635 94.285 ;
        RECT 63.815 93.725 64.645 94.045 ;
        RECT 63.405 93.210 63.665 93.530 ;
        RECT 63.815 93.355 64.530 93.725 ;
        RECT 64.300 93.070 64.530 93.355 ;
        RECT 64.785 93.530 65.015 94.285 ;
        RECT 65.195 93.725 66.025 94.045 ;
        RECT 64.785 93.210 65.045 93.530 ;
        RECT 65.195 93.355 65.910 93.725 ;
        RECT 65.680 93.070 65.910 93.355 ;
        RECT 66.165 93.530 66.395 94.285 ;
        RECT 66.575 93.725 67.405 94.045 ;
        RECT 66.165 93.210 66.425 93.530 ;
        RECT 66.575 93.355 67.290 93.725 ;
        RECT 67.060 93.070 67.290 93.355 ;
        RECT 67.545 93.530 67.775 94.285 ;
        RECT 67.955 93.725 68.785 94.045 ;
        RECT 67.545 93.210 67.805 93.530 ;
        RECT 67.955 93.070 68.670 93.725 ;
        RECT 68.925 93.530 69.155 94.285 ;
        RECT 68.925 93.210 69.185 93.530 ;
        RECT 37.525 92.770 37.825 92.880 ;
        RECT 40.090 92.770 40.350 92.845 ;
        RECT 37.525 92.600 40.350 92.770 ;
        RECT 37.525 92.490 37.825 92.600 ;
        RECT 40.090 92.525 40.350 92.600 ;
        RECT 55.535 92.840 56.735 93.070 ;
        RECT 57.400 92.840 58.115 93.070 ;
        RECT 58.780 92.840 59.495 93.070 ;
        RECT 60.160 92.840 60.875 93.070 ;
        RECT 61.540 92.840 62.255 93.070 ;
        RECT 62.920 92.840 63.635 93.070 ;
        RECT 64.300 92.840 65.015 93.070 ;
        RECT 65.680 92.840 66.395 93.070 ;
        RECT 67.060 92.840 67.775 93.070 ;
        RECT 36.025 92.350 36.325 92.460 ;
        RECT 44.590 92.350 44.850 92.425 ;
        RECT 36.025 92.180 44.850 92.350 ;
        RECT 36.025 92.070 36.325 92.180 ;
        RECT 44.590 92.105 44.850 92.180 ;
        RECT 55.535 92.005 56.225 92.840 ;
        RECT 38.590 91.995 38.850 92.005 ;
        RECT 38.590 91.930 39.370 91.995 ;
        RECT 43.090 91.930 43.350 92.005 ;
        RECT 37.590 91.760 43.350 91.930 ;
        RECT 55.905 91.820 56.365 91.865 ;
        RECT 38.590 91.695 39.370 91.760 ;
        RECT 38.590 91.685 38.850 91.695 ;
        RECT 43.090 91.685 43.350 91.760 ;
        RECT 55.535 91.590 56.365 91.820 ;
        RECT 31.545 91.035 31.805 91.110 ;
        RECT 35.560 91.035 35.880 91.080 ;
        RECT 31.545 90.865 35.880 91.035 ;
        RECT 31.545 90.790 31.805 90.865 ;
        RECT 35.560 90.820 35.880 90.865 ;
        RECT 36.045 91.035 36.305 91.110 ;
        RECT 37.090 91.035 37.350 91.110 ;
        RECT 36.045 90.865 37.350 91.035 ;
        RECT 36.045 90.790 36.305 90.865 ;
        RECT 37.090 90.790 37.350 90.865 ;
        RECT 39.045 91.035 39.305 91.110 ;
        RECT 40.545 91.035 40.805 91.110 ;
        RECT 42.025 91.035 42.325 91.145 ;
        RECT 39.045 90.865 42.325 91.035 ;
        RECT 39.045 90.790 39.305 90.865 ;
        RECT 40.545 90.790 40.805 90.865 ;
        RECT 42.025 90.755 42.325 90.865 ;
        RECT 43.545 91.035 43.805 91.110 ;
        RECT 45.045 91.035 45.305 91.110 ;
        RECT 46.525 91.035 46.825 91.145 ;
        RECT 47.785 91.035 48.085 91.145 ;
        RECT 43.545 90.865 48.085 91.035 ;
        RECT 43.545 90.790 43.805 90.865 ;
        RECT 45.045 90.790 45.305 90.865 ;
        RECT 46.525 90.755 46.825 90.865 ;
        RECT 47.785 90.755 48.085 90.865 ;
        RECT 47.155 90.405 47.455 90.515 ;
        RECT 49.675 90.405 49.975 90.515 ;
        RECT 47.155 90.235 49.975 90.405 ;
        RECT 47.155 90.125 47.455 90.235 ;
        RECT 49.675 90.125 49.975 90.235 ;
        RECT 47.785 89.775 48.085 89.885 ;
        RECT 50.305 89.775 50.605 89.885 ;
        RECT 47.785 89.605 50.605 89.775 ;
        RECT 47.785 89.495 48.085 89.605 ;
        RECT 50.305 89.495 50.605 89.605 ;
        RECT 33.085 89.230 33.345 89.305 ;
        RECT 34.090 89.230 34.350 89.305 ;
        RECT 33.085 89.060 34.350 89.230 ;
        RECT 33.085 88.985 33.345 89.060 ;
        RECT 34.090 88.985 34.350 89.060 ;
        RECT 35.275 88.100 35.575 88.490 ;
        RECT 38.275 88.100 38.575 88.490 ;
        RECT 41.275 88.100 41.575 88.490 ;
        RECT 44.275 88.100 44.575 88.490 ;
        RECT 42.025 87.810 42.325 87.920 ;
        RECT 47.155 87.810 47.455 87.920 ;
        RECT 42.025 87.640 47.455 87.810 ;
        RECT 54.450 87.750 55.200 88.440 ;
        RECT 55.535 87.755 55.765 91.590 ;
        RECT 55.905 91.545 56.365 91.590 ;
        RECT 55.905 89.885 56.365 89.930 ;
        RECT 56.505 89.885 56.735 92.840 ;
        RECT 56.915 92.005 57.605 92.700 ;
        RECT 57.285 91.820 57.745 91.865 ;
        RECT 55.905 89.655 56.735 89.885 ;
        RECT 56.915 91.590 57.745 91.820 ;
        RECT 55.905 89.610 56.365 89.655 ;
        RECT 42.025 87.530 42.325 87.640 ;
        RECT 47.155 87.530 47.455 87.640 ;
        RECT 33.775 87.050 34.075 87.440 ;
        RECT 36.775 87.050 37.075 87.440 ;
        RECT 39.775 87.050 40.075 87.440 ;
        RECT 42.775 87.050 43.075 87.440 ;
        RECT 45.775 87.050 46.075 87.440 ;
        RECT 54.480 86.940 55.170 87.750 ;
        RECT 55.535 87.105 55.855 87.755 ;
        RECT 56.045 86.940 56.735 89.465 ;
        RECT 56.915 87.755 57.145 91.590 ;
        RECT 57.285 91.545 57.745 91.590 ;
        RECT 57.285 89.885 57.745 89.930 ;
        RECT 57.885 89.885 58.115 92.840 ;
        RECT 58.295 92.005 58.985 92.700 ;
        RECT 58.665 91.820 59.125 91.865 ;
        RECT 57.285 89.655 58.115 89.885 ;
        RECT 58.295 91.590 59.125 91.820 ;
        RECT 57.285 89.610 57.745 89.655 ;
        RECT 57.425 88.775 58.115 89.465 ;
        RECT 57.425 87.915 58.115 88.605 ;
        RECT 58.295 87.755 58.525 91.590 ;
        RECT 58.665 91.545 59.125 91.590 ;
        RECT 58.665 89.885 59.125 89.930 ;
        RECT 59.265 89.885 59.495 92.840 ;
        RECT 59.675 92.005 60.365 92.700 ;
        RECT 60.045 91.820 60.505 91.865 ;
        RECT 58.665 89.655 59.495 89.885 ;
        RECT 59.675 91.590 60.505 91.820 ;
        RECT 58.665 89.610 59.125 89.655 ;
        RECT 58.805 88.775 59.495 89.465 ;
        RECT 58.805 87.915 59.495 88.605 ;
        RECT 59.675 87.755 59.905 91.590 ;
        RECT 60.045 91.545 60.505 91.590 ;
        RECT 60.045 89.885 60.505 89.930 ;
        RECT 60.645 89.885 60.875 92.840 ;
        RECT 61.055 92.005 61.745 92.700 ;
        RECT 61.425 91.820 61.885 91.865 ;
        RECT 60.045 89.655 60.875 89.885 ;
        RECT 61.055 91.590 61.885 91.820 ;
        RECT 60.045 89.610 60.505 89.655 ;
        RECT 60.185 88.775 60.875 89.465 ;
        RECT 60.185 87.915 60.875 88.605 ;
        RECT 61.055 87.755 61.285 91.590 ;
        RECT 61.425 91.545 61.885 91.590 ;
        RECT 61.425 89.885 61.885 89.930 ;
        RECT 62.025 89.885 62.255 92.840 ;
        RECT 62.435 92.005 63.125 92.700 ;
        RECT 62.805 91.820 63.265 91.865 ;
        RECT 61.425 89.655 62.255 89.885 ;
        RECT 62.435 91.590 63.265 91.820 ;
        RECT 61.425 89.610 61.885 89.655 ;
        RECT 61.565 88.775 62.255 89.465 ;
        RECT 61.565 87.915 62.255 88.605 ;
        RECT 62.435 87.755 62.665 91.590 ;
        RECT 62.805 91.545 63.265 91.590 ;
        RECT 62.805 89.885 63.265 89.930 ;
        RECT 63.405 89.885 63.635 92.840 ;
        RECT 63.815 92.005 64.505 92.700 ;
        RECT 64.185 91.820 64.645 91.865 ;
        RECT 62.805 89.655 63.635 89.885 ;
        RECT 63.815 91.590 64.645 91.820 ;
        RECT 62.805 89.610 63.265 89.655 ;
        RECT 62.945 88.775 63.635 89.465 ;
        RECT 62.945 87.915 63.635 88.605 ;
        RECT 63.815 87.755 64.045 91.590 ;
        RECT 64.185 91.545 64.645 91.590 ;
        RECT 64.185 89.885 64.645 89.930 ;
        RECT 64.785 89.885 65.015 92.840 ;
        RECT 65.195 92.005 65.885 92.700 ;
        RECT 65.565 91.820 66.025 91.865 ;
        RECT 64.185 89.655 65.015 89.885 ;
        RECT 65.195 91.590 66.025 91.820 ;
        RECT 64.185 89.610 64.645 89.655 ;
        RECT 64.325 88.775 65.015 89.465 ;
        RECT 64.325 87.915 65.015 88.605 ;
        RECT 65.195 87.755 65.425 91.590 ;
        RECT 65.565 91.545 66.025 91.590 ;
        RECT 65.565 89.885 66.025 89.930 ;
        RECT 66.165 89.885 66.395 92.840 ;
        RECT 66.575 92.005 67.265 92.700 ;
        RECT 66.945 91.820 67.405 91.865 ;
        RECT 65.565 89.655 66.395 89.885 ;
        RECT 66.575 91.590 67.405 91.820 ;
        RECT 65.565 89.610 66.025 89.655 ;
        RECT 65.705 88.775 66.395 89.465 ;
        RECT 65.705 87.915 66.395 88.605 ;
        RECT 66.575 87.755 66.805 91.590 ;
        RECT 66.945 91.545 67.405 91.590 ;
        RECT 66.945 89.885 67.405 89.930 ;
        RECT 67.545 89.885 67.775 92.840 ;
        RECT 67.955 92.840 69.155 93.070 ;
        RECT 67.955 92.005 68.645 92.840 ;
        RECT 68.325 91.820 68.785 91.865 ;
        RECT 66.945 89.655 67.775 89.885 ;
        RECT 67.955 91.590 68.785 91.820 ;
        RECT 66.945 89.610 67.405 89.655 ;
        RECT 67.085 88.775 67.775 89.465 ;
        RECT 67.085 87.915 67.775 88.605 ;
        RECT 67.955 87.755 68.185 91.590 ;
        RECT 68.325 91.545 68.785 91.590 ;
        RECT 68.325 89.885 68.785 89.930 ;
        RECT 68.925 89.885 69.155 92.840 ;
        RECT 68.325 89.655 69.155 89.885 ;
        RECT 68.325 89.610 68.785 89.655 ;
        RECT 56.915 87.105 57.235 87.755 ;
        RECT 58.295 87.105 58.615 87.755 ;
        RECT 59.675 87.105 59.995 87.755 ;
        RECT 61.055 87.105 61.375 87.755 ;
        RECT 62.435 87.105 62.755 87.755 ;
        RECT 63.815 87.105 64.135 87.755 ;
        RECT 65.195 87.105 65.515 87.755 ;
        RECT 66.575 87.105 66.895 87.755 ;
        RECT 67.955 87.105 68.275 87.755 ;
        RECT 68.465 86.940 69.155 89.465 ;
        RECT 70.655 86.940 71.345 86.985 ;
        RECT 34.525 86.480 34.825 86.590 ;
        RECT 41.590 86.480 41.850 86.555 ;
        RECT 46.090 86.480 46.350 86.555 ;
        RECT 34.525 86.310 46.350 86.480 ;
        RECT 34.525 86.200 34.825 86.310 ;
        RECT 41.590 86.235 41.850 86.310 ;
        RECT 46.090 86.235 46.350 86.310 ;
        RECT 54.480 86.250 71.345 86.940 ;
        RECT 70.655 86.205 71.345 86.250 ;
        RECT 37.525 86.060 37.825 86.170 ;
        RECT 40.090 86.060 40.350 86.135 ;
        RECT 37.525 85.890 40.350 86.060 ;
        RECT 37.525 85.780 37.825 85.890 ;
        RECT 40.090 85.815 40.350 85.890 ;
        RECT 36.025 85.640 36.325 85.750 ;
        RECT 50.600 85.740 50.900 85.785 ;
        RECT 52.260 85.740 52.560 85.785 ;
        RECT 53.920 85.740 54.220 85.785 ;
        RECT 55.580 85.740 55.880 85.785 ;
        RECT 57.240 85.740 57.540 85.785 ;
        RECT 58.900 85.740 59.200 85.785 ;
        RECT 44.590 85.640 44.850 85.715 ;
        RECT 36.025 85.470 44.850 85.640 ;
        RECT 36.025 85.360 36.325 85.470 ;
        RECT 44.590 85.395 44.850 85.470 ;
        RECT 50.570 85.440 50.930 85.740 ;
        RECT 52.230 85.440 52.590 85.740 ;
        RECT 53.890 85.440 54.250 85.740 ;
        RECT 55.550 85.440 55.910 85.740 ;
        RECT 57.210 85.440 57.570 85.740 ;
        RECT 58.870 85.440 59.230 85.740 ;
        RECT 50.600 85.395 50.900 85.440 ;
        RECT 52.260 85.395 52.560 85.440 ;
        RECT 53.920 85.395 54.220 85.440 ;
        RECT 55.580 85.395 55.880 85.440 ;
        RECT 57.240 85.395 57.540 85.440 ;
        RECT 58.900 85.395 59.200 85.440 ;
        RECT 60.560 85.325 60.860 85.370 ;
        RECT 36.450 85.220 36.710 85.290 ;
        RECT 38.590 85.220 38.850 85.295 ;
        RECT 43.090 85.220 43.350 85.295 ;
        RECT 36.090 85.050 43.350 85.220 ;
        RECT 36.450 84.970 36.710 85.050 ;
        RECT 38.590 84.975 38.850 85.050 ;
        RECT 43.090 84.975 43.350 85.050 ;
        RECT 60.530 85.025 60.890 85.325 ;
        RECT 60.560 84.980 60.860 85.025 ;
        RECT 62.220 84.700 62.520 84.745 ;
        RECT 31.930 84.325 32.190 84.400 ;
        RECT 35.560 84.325 35.880 84.370 ;
        RECT 31.930 84.155 35.880 84.325 ;
        RECT 31.930 84.080 32.190 84.155 ;
        RECT 35.560 84.110 35.880 84.155 ;
        RECT 36.045 84.325 36.305 84.400 ;
        RECT 37.090 84.325 37.350 84.400 ;
        RECT 36.045 84.155 37.350 84.325 ;
        RECT 36.045 84.080 36.305 84.155 ;
        RECT 37.090 84.080 37.350 84.155 ;
        RECT 39.045 84.325 39.305 84.400 ;
        RECT 40.545 84.325 40.805 84.400 ;
        RECT 42.025 84.325 42.325 84.435 ;
        RECT 39.045 84.155 42.325 84.325 ;
        RECT 39.045 84.080 39.305 84.155 ;
        RECT 40.545 84.080 40.805 84.155 ;
        RECT 42.025 84.045 42.325 84.155 ;
        RECT 43.545 84.325 43.805 84.400 ;
        RECT 45.045 84.325 45.305 84.400 ;
        RECT 46.525 84.325 46.825 84.435 ;
        RECT 47.785 84.325 48.085 84.435 ;
        RECT 62.190 84.400 62.550 84.700 ;
        RECT 62.220 84.355 62.520 84.400 ;
        RECT 43.545 84.155 48.085 84.325 ;
        RECT 43.545 84.080 43.805 84.155 ;
        RECT 45.045 84.080 45.305 84.155 ;
        RECT 46.525 84.045 46.825 84.155 ;
        RECT 47.785 84.045 48.085 84.155 ;
        RECT 37.545 82.520 37.805 82.595 ;
        RECT 39.025 82.520 39.325 82.630 ;
        RECT 37.545 82.350 39.325 82.520 ;
        RECT 37.545 82.275 37.805 82.350 ;
        RECT 39.025 82.240 39.325 82.350 ;
        RECT 35.275 81.390 35.575 81.780 ;
        RECT 38.275 81.390 38.575 81.780 ;
        RECT 41.275 81.390 41.575 81.780 ;
        RECT 44.275 81.390 44.575 81.780 ;
        RECT 42.025 81.100 42.325 81.210 ;
        RECT 48.415 81.100 48.715 81.210 ;
        RECT 42.025 80.930 48.715 81.100 ;
        RECT 42.025 80.820 42.325 80.930 ;
        RECT 48.415 80.820 48.715 80.930 ;
        RECT 33.775 80.340 34.075 80.730 ;
        RECT 36.775 80.340 37.075 80.730 ;
        RECT 39.775 80.340 40.075 80.730 ;
        RECT 42.775 80.340 43.075 80.730 ;
        RECT 45.775 80.340 46.075 80.730 ;
        RECT 34.525 79.770 34.825 79.880 ;
        RECT 41.590 79.770 41.850 79.845 ;
        RECT 46.090 79.770 46.350 79.845 ;
        RECT 34.525 79.600 46.350 79.770 ;
        RECT 34.525 79.490 34.825 79.600 ;
        RECT 41.590 79.525 41.850 79.600 ;
        RECT 46.090 79.525 46.350 79.600 ;
        RECT 37.525 79.350 37.825 79.460 ;
        RECT 40.090 79.350 40.350 79.425 ;
        RECT 37.525 79.180 40.350 79.350 ;
        RECT 37.525 79.070 37.825 79.180 ;
        RECT 40.090 79.105 40.350 79.180 ;
        RECT 36.025 78.930 36.325 79.040 ;
        RECT 44.590 78.930 44.850 79.005 ;
        RECT 36.025 78.760 44.850 78.930 ;
        RECT 36.025 78.650 36.325 78.760 ;
        RECT 44.590 78.685 44.850 78.760 ;
        RECT 38.590 78.575 38.850 78.585 ;
        RECT 38.590 78.510 39.370 78.575 ;
        RECT 43.090 78.510 43.350 78.585 ;
        RECT 37.590 78.340 43.350 78.510 ;
        RECT 38.590 78.275 39.370 78.340 ;
        RECT 38.590 78.265 38.850 78.275 ;
        RECT 43.090 78.265 43.350 78.340 ;
        RECT 31.545 77.615 31.805 77.690 ;
        RECT 35.560 77.615 35.880 77.660 ;
        RECT 31.545 77.445 35.880 77.615 ;
        RECT 31.545 77.370 31.805 77.445 ;
        RECT 35.560 77.400 35.880 77.445 ;
        RECT 36.045 77.615 36.305 77.690 ;
        RECT 37.090 77.615 37.350 77.690 ;
        RECT 36.045 77.445 37.350 77.615 ;
        RECT 36.045 77.370 36.305 77.445 ;
        RECT 37.090 77.370 37.350 77.445 ;
        RECT 39.045 77.615 39.305 77.690 ;
        RECT 40.545 77.615 40.805 77.690 ;
        RECT 42.025 77.615 42.325 77.725 ;
        RECT 39.045 77.445 42.325 77.615 ;
        RECT 39.045 77.370 39.305 77.445 ;
        RECT 40.545 77.370 40.805 77.445 ;
        RECT 42.025 77.335 42.325 77.445 ;
        RECT 43.545 77.615 43.805 77.690 ;
        RECT 45.045 77.615 45.305 77.690 ;
        RECT 46.525 77.615 46.825 77.725 ;
        RECT 49.045 77.615 49.345 77.725 ;
        RECT 43.545 77.445 49.345 77.615 ;
        RECT 43.545 77.370 43.805 77.445 ;
        RECT 45.045 77.370 45.305 77.445 ;
        RECT 46.525 77.335 46.825 77.445 ;
        RECT 49.045 77.335 49.345 77.445 ;
        RECT 32.700 75.810 32.960 75.885 ;
        RECT 34.090 75.810 34.350 75.885 ;
        RECT 32.700 75.640 34.350 75.810 ;
        RECT 32.700 75.565 32.960 75.640 ;
        RECT 34.090 75.565 34.350 75.640 ;
        RECT 35.275 74.680 35.575 75.070 ;
        RECT 38.275 74.680 38.575 75.070 ;
        RECT 41.275 74.680 41.575 75.070 ;
        RECT 44.275 74.680 44.575 75.070 ;
        RECT 42.025 74.390 42.325 74.500 ;
        RECT 51.565 74.390 51.865 74.500 ;
        RECT 42.025 74.220 51.865 74.390 ;
        RECT 42.025 74.110 42.325 74.220 ;
        RECT 51.565 74.110 51.865 74.220 ;
        RECT 33.775 73.630 34.075 74.020 ;
        RECT 36.775 73.630 37.075 74.020 ;
        RECT 39.775 73.630 40.075 74.020 ;
        RECT 42.775 73.630 43.075 74.020 ;
        RECT 45.775 73.630 46.075 74.020 ;
        RECT 34.525 73.060 34.825 73.170 ;
        RECT 41.590 73.060 41.850 73.135 ;
        RECT 46.090 73.060 46.350 73.135 ;
        RECT 34.525 72.890 46.350 73.060 ;
        RECT 34.525 72.780 34.825 72.890 ;
        RECT 41.590 72.815 41.850 72.890 ;
        RECT 46.090 72.815 46.350 72.890 ;
        RECT 37.525 72.640 37.825 72.750 ;
        RECT 40.090 72.640 40.350 72.715 ;
        RECT 37.525 72.470 40.350 72.640 ;
        RECT 37.525 72.360 37.825 72.470 ;
        RECT 40.090 72.395 40.350 72.470 ;
        RECT 36.025 72.220 36.325 72.330 ;
        RECT 44.590 72.220 44.850 72.295 ;
        RECT 36.025 72.050 44.850 72.220 ;
        RECT 36.025 71.940 36.325 72.050 ;
        RECT 44.590 71.975 44.850 72.050 ;
        RECT 36.450 71.800 36.710 71.870 ;
        RECT 38.590 71.800 38.850 71.875 ;
        RECT 43.090 71.800 43.350 71.875 ;
        RECT 36.090 71.630 43.350 71.800 ;
        RECT 36.450 71.550 36.710 71.630 ;
        RECT 38.590 71.555 38.850 71.630 ;
        RECT 43.090 71.555 43.350 71.630 ;
        RECT 31.900 70.905 32.220 70.950 ;
        RECT 35.560 70.905 35.880 70.950 ;
        RECT 31.900 70.735 35.880 70.905 ;
        RECT 31.900 70.690 32.220 70.735 ;
        RECT 35.560 70.690 35.880 70.735 ;
        RECT 36.045 70.905 36.305 70.980 ;
        RECT 37.090 70.905 37.350 70.980 ;
        RECT 36.045 70.735 37.350 70.905 ;
        RECT 36.045 70.660 36.305 70.735 ;
        RECT 37.090 70.660 37.350 70.735 ;
        RECT 39.045 70.905 39.305 70.980 ;
        RECT 40.545 70.905 40.805 70.980 ;
        RECT 42.025 70.905 42.325 71.015 ;
        RECT 39.045 70.735 42.325 70.905 ;
        RECT 39.045 70.660 39.305 70.735 ;
        RECT 40.545 70.660 40.805 70.735 ;
        RECT 42.025 70.625 42.325 70.735 ;
        RECT 43.545 70.905 43.805 70.980 ;
        RECT 45.045 70.905 45.305 70.980 ;
        RECT 46.525 70.905 46.825 71.015 ;
        RECT 50.935 70.905 51.235 71.015 ;
        RECT 43.545 70.735 51.235 70.905 ;
        RECT 43.545 70.660 43.805 70.735 ;
        RECT 45.045 70.660 45.305 70.735 ;
        RECT 46.525 70.625 46.825 70.735 ;
        RECT 50.935 70.625 51.235 70.735 ;
        RECT 37.545 69.100 37.805 69.175 ;
        RECT 39.025 69.100 39.325 69.210 ;
        RECT 37.545 68.930 39.325 69.100 ;
        RECT 37.545 68.855 37.805 68.930 ;
        RECT 39.025 68.820 39.325 68.930 ;
        RECT 35.275 67.970 35.575 68.360 ;
        RECT 38.275 67.970 38.575 68.360 ;
        RECT 41.275 67.970 41.575 68.360 ;
        RECT 44.275 67.970 44.575 68.360 ;
        RECT 42.025 67.680 42.325 67.790 ;
        RECT 47.155 67.680 47.455 67.790 ;
        RECT 42.025 67.510 47.455 67.680 ;
        RECT 42.025 67.400 42.325 67.510 ;
        RECT 47.155 67.400 47.455 67.510 ;
        RECT 33.775 66.920 34.075 67.310 ;
        RECT 36.775 66.920 37.075 67.310 ;
        RECT 39.775 66.920 40.075 67.310 ;
        RECT 42.775 66.920 43.075 67.310 ;
        RECT 45.775 66.920 46.075 67.310 ;
        RECT 34.525 66.350 34.825 66.460 ;
        RECT 41.590 66.350 41.850 66.425 ;
        RECT 46.090 66.350 46.350 66.425 ;
        RECT 34.525 66.180 46.350 66.350 ;
        RECT 34.525 66.070 34.825 66.180 ;
        RECT 41.590 66.105 41.850 66.180 ;
        RECT 46.090 66.105 46.350 66.180 ;
        RECT 37.525 65.930 37.825 66.040 ;
        RECT 40.090 65.930 40.350 66.005 ;
        RECT 37.525 65.760 40.350 65.930 ;
        RECT 37.525 65.650 37.825 65.760 ;
        RECT 40.090 65.685 40.350 65.760 ;
        RECT 36.025 65.510 36.325 65.620 ;
        RECT 44.590 65.510 44.850 65.585 ;
        RECT 36.025 65.340 44.850 65.510 ;
        RECT 36.025 65.230 36.325 65.340 ;
        RECT 44.590 65.265 44.850 65.340 ;
        RECT 38.590 65.155 38.850 65.165 ;
        RECT 38.590 65.090 39.370 65.155 ;
        RECT 43.090 65.090 43.350 65.165 ;
        RECT 37.590 64.920 43.350 65.090 ;
        RECT 38.590 64.855 39.370 64.920 ;
        RECT 38.590 64.845 38.850 64.855 ;
        RECT 43.090 64.845 43.350 64.920 ;
        RECT 31.545 64.195 31.805 64.270 ;
        RECT 35.560 64.195 35.880 64.240 ;
        RECT 31.545 64.025 35.880 64.195 ;
        RECT 31.545 63.950 31.805 64.025 ;
        RECT 35.560 63.980 35.880 64.025 ;
        RECT 36.045 64.195 36.305 64.270 ;
        RECT 37.090 64.195 37.350 64.270 ;
        RECT 36.045 64.025 37.350 64.195 ;
        RECT 36.045 63.950 36.305 64.025 ;
        RECT 37.090 63.950 37.350 64.025 ;
        RECT 39.045 64.195 39.305 64.270 ;
        RECT 40.545 64.195 40.805 64.270 ;
        RECT 42.025 64.195 42.325 64.305 ;
        RECT 39.045 64.025 42.325 64.195 ;
        RECT 39.045 63.950 39.305 64.025 ;
        RECT 40.545 63.950 40.805 64.025 ;
        RECT 42.025 63.915 42.325 64.025 ;
        RECT 43.545 64.195 43.805 64.270 ;
        RECT 45.045 64.195 45.305 64.270 ;
        RECT 46.525 64.195 46.825 64.305 ;
        RECT 47.785 64.195 48.085 64.305 ;
        RECT 43.545 64.025 48.085 64.195 ;
        RECT 43.545 63.950 43.805 64.025 ;
        RECT 45.045 63.950 45.305 64.025 ;
        RECT 46.525 63.915 46.825 64.025 ;
        RECT 47.785 63.915 48.085 64.025 ;
        RECT 32.315 62.390 32.575 62.465 ;
        RECT 34.090 62.390 34.350 62.465 ;
        RECT 32.315 62.220 34.350 62.390 ;
        RECT 32.315 62.145 32.575 62.220 ;
        RECT 34.090 62.145 34.350 62.220 ;
        RECT 35.275 61.260 35.575 61.650 ;
        RECT 38.275 61.260 38.575 61.650 ;
        RECT 41.275 61.260 41.575 61.650 ;
        RECT 44.275 61.260 44.575 61.650 ;
        RECT 42.025 60.970 42.325 61.080 ;
        RECT 49.045 60.970 49.345 61.080 ;
        RECT 42.025 60.800 49.345 60.970 ;
        RECT 42.025 60.690 42.325 60.800 ;
        RECT 49.045 60.690 49.345 60.800 ;
        RECT 33.775 60.210 34.075 60.600 ;
        RECT 36.775 60.210 37.075 60.600 ;
        RECT 39.775 60.210 40.075 60.600 ;
        RECT 42.775 60.210 43.075 60.600 ;
        RECT 45.775 60.210 46.075 60.600 ;
        RECT 34.525 59.640 34.825 59.750 ;
        RECT 41.590 59.640 41.850 59.715 ;
        RECT 46.090 59.640 46.350 59.715 ;
        RECT 34.525 59.470 46.350 59.640 ;
        RECT 34.525 59.360 34.825 59.470 ;
        RECT 41.590 59.395 41.850 59.470 ;
        RECT 46.090 59.395 46.350 59.470 ;
        RECT 37.525 59.220 37.825 59.330 ;
        RECT 40.090 59.220 40.350 59.295 ;
        RECT 37.525 59.050 40.350 59.220 ;
        RECT 37.525 58.940 37.825 59.050 ;
        RECT 40.090 58.975 40.350 59.050 ;
        RECT 36.025 58.800 36.325 58.910 ;
        RECT 44.590 58.800 44.850 58.875 ;
        RECT 36.025 58.630 44.850 58.800 ;
        RECT 36.025 58.520 36.325 58.630 ;
        RECT 44.590 58.555 44.850 58.630 ;
        RECT 36.450 58.380 36.710 58.450 ;
        RECT 38.590 58.380 38.850 58.455 ;
        RECT 43.090 58.380 43.350 58.455 ;
        RECT 36.090 58.210 43.350 58.380 ;
        RECT 36.450 58.130 36.710 58.210 ;
        RECT 38.590 58.135 38.850 58.210 ;
        RECT 43.090 58.135 43.350 58.210 ;
        RECT 28.645 57.485 28.965 57.530 ;
        RECT 31.930 57.485 32.190 57.560 ;
        RECT 35.560 57.485 35.880 57.530 ;
        RECT 28.645 57.315 35.880 57.485 ;
        RECT 28.645 57.270 28.965 57.315 ;
        RECT 31.930 57.240 32.190 57.315 ;
        RECT 35.560 57.270 35.880 57.315 ;
        RECT 36.045 57.485 36.305 57.560 ;
        RECT 37.090 57.485 37.350 57.560 ;
        RECT 36.045 57.315 37.350 57.485 ;
        RECT 36.045 57.240 36.305 57.315 ;
        RECT 37.090 57.240 37.350 57.315 ;
        RECT 39.045 57.485 39.305 57.560 ;
        RECT 40.545 57.485 40.805 57.560 ;
        RECT 42.025 57.485 42.325 57.595 ;
        RECT 39.045 57.315 42.325 57.485 ;
        RECT 39.045 57.240 39.305 57.315 ;
        RECT 40.545 57.240 40.805 57.315 ;
        RECT 42.025 57.205 42.325 57.315 ;
        RECT 43.545 57.485 43.805 57.560 ;
        RECT 45.045 57.485 45.305 57.560 ;
        RECT 46.525 57.485 46.825 57.595 ;
        RECT 48.415 57.485 48.715 57.595 ;
        RECT 43.545 57.315 48.715 57.485 ;
        RECT 43.545 57.240 43.805 57.315 ;
        RECT 45.045 57.240 45.305 57.315 ;
        RECT 46.525 57.205 46.825 57.315 ;
        RECT 48.415 57.205 48.715 57.315 ;
        RECT 37.545 55.680 37.805 55.755 ;
        RECT 39.025 55.680 39.325 55.790 ;
        RECT 37.545 55.510 39.325 55.680 ;
        RECT 37.545 55.435 37.805 55.510 ;
        RECT 39.025 55.400 39.325 55.510 ;
        RECT 35.275 54.550 35.575 54.940 ;
        RECT 38.275 54.550 38.575 54.940 ;
        RECT 41.275 54.550 41.575 54.940 ;
        RECT 44.275 54.550 44.575 54.940 ;
        RECT 42.025 54.260 42.325 54.370 ;
        RECT 50.305 54.260 50.605 54.370 ;
        RECT 42.025 54.090 50.605 54.260 ;
        RECT 42.025 53.980 42.325 54.090 ;
        RECT 50.305 53.980 50.605 54.090 ;
        RECT 33.775 53.500 34.075 53.890 ;
        RECT 36.775 53.500 37.075 53.890 ;
        RECT 39.775 53.500 40.075 53.890 ;
        RECT 42.775 53.500 43.075 53.890 ;
        RECT 45.775 53.500 46.075 53.890 ;
        RECT 63.050 53.130 63.350 53.175 ;
        RECT 34.525 52.930 34.825 53.040 ;
        RECT 41.590 52.930 41.850 53.005 ;
        RECT 46.090 52.930 46.350 53.005 ;
        RECT 34.525 52.760 46.350 52.930 ;
        RECT 63.020 52.830 63.380 53.130 ;
        RECT 63.050 52.785 63.350 52.830 ;
        RECT 34.525 52.650 34.825 52.760 ;
        RECT 41.590 52.685 41.850 52.760 ;
        RECT 46.090 52.685 46.350 52.760 ;
        RECT 37.525 52.510 37.825 52.620 ;
        RECT 40.090 52.510 40.350 52.585 ;
        RECT 37.525 52.340 40.350 52.510 ;
        RECT 61.390 52.505 61.690 52.550 ;
        RECT 37.525 52.230 37.825 52.340 ;
        RECT 40.090 52.265 40.350 52.340 ;
        RECT 61.360 52.205 61.720 52.505 ;
        RECT 36.025 52.090 36.325 52.200 ;
        RECT 44.590 52.090 44.850 52.165 ;
        RECT 61.390 52.160 61.690 52.205 ;
        RECT 36.025 51.920 44.850 52.090 ;
        RECT 36.025 51.810 36.325 51.920 ;
        RECT 44.590 51.845 44.850 51.920 ;
        RECT 59.730 51.880 60.030 51.925 ;
        RECT 38.590 51.735 38.850 51.745 ;
        RECT 38.590 51.670 39.370 51.735 ;
        RECT 43.090 51.670 43.350 51.745 ;
        RECT 37.590 51.500 43.350 51.670 ;
        RECT 59.700 51.580 60.060 51.880 ;
        RECT 59.730 51.535 60.030 51.580 ;
        RECT 38.590 51.435 39.370 51.500 ;
        RECT 38.590 51.425 38.850 51.435 ;
        RECT 43.090 51.425 43.350 51.500 ;
        RECT 58.070 50.910 58.370 51.300 ;
        RECT 28.645 50.775 28.965 50.820 ;
        RECT 31.545 50.775 31.805 50.850 ;
        RECT 35.560 50.775 35.880 50.820 ;
        RECT 28.645 50.605 35.880 50.775 ;
        RECT 28.645 50.560 28.965 50.605 ;
        RECT 31.545 50.530 31.805 50.605 ;
        RECT 35.560 50.560 35.880 50.605 ;
        RECT 36.045 50.775 36.305 50.850 ;
        RECT 37.090 50.775 37.350 50.850 ;
        RECT 36.045 50.605 37.350 50.775 ;
        RECT 36.045 50.530 36.305 50.605 ;
        RECT 37.090 50.530 37.350 50.605 ;
        RECT 39.045 50.775 39.305 50.850 ;
        RECT 40.545 50.775 40.805 50.850 ;
        RECT 42.025 50.775 42.325 50.885 ;
        RECT 39.045 50.605 42.325 50.775 ;
        RECT 39.045 50.530 39.305 50.605 ;
        RECT 40.545 50.530 40.805 50.605 ;
        RECT 42.025 50.495 42.325 50.605 ;
        RECT 43.545 50.775 43.805 50.850 ;
        RECT 45.045 50.775 45.305 50.850 ;
        RECT 46.525 50.775 46.825 50.885 ;
        RECT 49.675 50.775 49.975 50.885 ;
        RECT 43.545 50.605 49.975 50.775 ;
        RECT 43.545 50.530 43.805 50.605 ;
        RECT 45.045 50.530 45.305 50.605 ;
        RECT 46.525 50.495 46.825 50.605 ;
        RECT 49.675 50.495 49.975 50.605 ;
        RECT 51.305 50.385 55.955 50.885 ;
        RECT 56.410 50.630 56.710 50.675 ;
        RECT 31.930 48.970 32.190 49.045 ;
        RECT 34.090 48.970 34.350 49.045 ;
        RECT 31.930 48.800 34.350 48.970 ;
        RECT 51.305 48.865 51.805 50.385 ;
        RECT 55.455 50.080 55.955 50.385 ;
        RECT 56.380 50.330 56.740 50.630 ;
        RECT 56.410 50.285 56.710 50.330 ;
        RECT 62.170 50.080 62.670 50.110 ;
        RECT 54.750 50.005 55.050 50.050 ;
        RECT 54.720 49.705 55.080 50.005 ;
        RECT 54.750 49.660 55.050 49.705 ;
        RECT 55.455 49.580 62.670 50.080 ;
        RECT 62.170 49.550 62.670 49.580 ;
        RECT 53.090 49.380 53.390 49.425 ;
        RECT 53.060 49.080 53.420 49.380 ;
        RECT 53.090 49.035 53.390 49.080 ;
        RECT 65.655 49.025 66.345 54.890 ;
        RECT 68.810 49.820 69.160 51.740 ;
        RECT 68.810 49.580 69.935 49.820 ;
        RECT 31.930 48.725 32.190 48.800 ;
        RECT 34.090 48.725 34.350 48.800 ;
        RECT 49.330 48.365 51.805 48.865 ;
        RECT 53.720 48.755 54.020 48.800 ;
        RECT 53.690 48.455 54.050 48.755 ;
        RECT 53.720 48.410 54.020 48.455 ;
        RECT 35.275 47.840 35.575 48.230 ;
        RECT 38.275 47.840 38.575 48.230 ;
        RECT 41.275 47.840 41.575 48.230 ;
        RECT 44.275 47.840 44.575 48.230 ;
        RECT 32.700 47.550 32.960 47.625 ;
        RECT 42.025 47.550 42.325 47.660 ;
        RECT 32.700 47.380 42.325 47.550 ;
        RECT 32.700 47.305 32.960 47.380 ;
        RECT 42.025 47.270 42.325 47.380 ;
        RECT 33.775 46.790 34.075 47.180 ;
        RECT 36.775 46.790 37.075 47.180 ;
        RECT 39.775 46.790 40.075 47.180 ;
        RECT 42.775 46.790 43.075 47.180 ;
        RECT 45.775 46.790 46.075 47.180 ;
        RECT 34.525 46.220 34.825 46.330 ;
        RECT 41.590 46.220 41.850 46.295 ;
        RECT 46.090 46.220 46.350 46.295 ;
        RECT 34.525 46.050 46.350 46.220 ;
        RECT 34.525 45.940 34.825 46.050 ;
        RECT 41.590 45.975 41.850 46.050 ;
        RECT 46.090 45.975 46.350 46.050 ;
        RECT 37.525 45.800 37.825 45.910 ;
        RECT 40.090 45.800 40.350 45.875 ;
        RECT 37.525 45.630 40.350 45.800 ;
        RECT 37.525 45.520 37.825 45.630 ;
        RECT 40.090 45.555 40.350 45.630 ;
        RECT 36.025 45.380 36.325 45.490 ;
        RECT 44.590 45.380 44.850 45.455 ;
        RECT 36.025 45.210 44.850 45.380 ;
        RECT 36.025 45.100 36.325 45.210 ;
        RECT 44.590 45.135 44.850 45.210 ;
        RECT 36.450 44.960 36.710 45.030 ;
        RECT 38.590 44.960 38.850 45.035 ;
        RECT 43.090 44.960 43.350 45.035 ;
        RECT 36.090 44.790 43.350 44.960 ;
        RECT 36.450 44.710 36.710 44.790 ;
        RECT 38.590 44.715 38.850 44.790 ;
        RECT 43.090 44.715 43.350 44.790 ;
        RECT 33.085 44.485 33.345 44.560 ;
        RECT 33.085 44.315 43.760 44.485 ;
        RECT 33.085 44.240 33.345 44.315 ;
        RECT 20.480 43.805 20.890 44.155 ;
        RECT 28.645 44.065 28.965 44.110 ;
        RECT 35.560 44.065 35.880 44.110 ;
        RECT 28.645 43.895 35.880 44.065 ;
        RECT 28.645 43.850 28.965 43.895 ;
        RECT 35.560 43.850 35.880 43.895 ;
        RECT 36.045 44.065 36.305 44.140 ;
        RECT 37.090 44.065 37.350 44.140 ;
        RECT 36.045 43.895 37.350 44.065 ;
        RECT 36.045 43.820 36.305 43.895 ;
        RECT 37.090 43.820 37.350 43.895 ;
        RECT 39.045 44.065 39.305 44.140 ;
        RECT 40.545 44.065 40.805 44.140 ;
        RECT 42.025 44.065 42.325 44.175 ;
        RECT 43.590 44.140 43.760 44.315 ;
        RECT 39.045 43.895 42.325 44.065 ;
        RECT 39.045 43.820 39.305 43.895 ;
        RECT 40.545 43.820 40.805 43.895 ;
        RECT 42.025 43.785 42.325 43.895 ;
        RECT 43.545 44.065 43.805 44.140 ;
        RECT 45.045 44.065 45.305 44.140 ;
        RECT 46.525 44.065 46.825 44.175 ;
        RECT 43.545 43.895 46.825 44.065 ;
        RECT 43.545 43.820 43.805 43.895 ;
        RECT 45.045 43.820 45.305 43.895 ;
        RECT 46.525 43.785 46.825 43.895 ;
        RECT 37.545 42.260 37.805 42.335 ;
        RECT 39.025 42.260 39.325 42.370 ;
        RECT 37.545 42.090 39.325 42.260 ;
        RECT 37.545 42.015 37.805 42.090 ;
        RECT 39.025 41.980 39.325 42.090 ;
        RECT 35.275 41.130 35.575 41.520 ;
        RECT 38.275 41.130 38.575 41.520 ;
        RECT 41.275 41.130 41.575 41.520 ;
        RECT 44.275 41.130 44.575 41.520 ;
        RECT 31.930 40.840 32.190 40.915 ;
        RECT 42.025 40.840 42.325 40.950 ;
        RECT 31.930 40.670 42.325 40.840 ;
        RECT 31.930 40.595 32.190 40.670 ;
        RECT 42.025 40.560 42.325 40.670 ;
        RECT 33.775 40.080 34.075 40.470 ;
        RECT 36.775 40.080 37.075 40.470 ;
        RECT 39.775 40.080 40.075 40.470 ;
        RECT 42.775 40.080 43.075 40.470 ;
        RECT 45.775 40.080 46.075 40.470 ;
        RECT 34.525 39.510 34.825 39.620 ;
        RECT 41.590 39.510 41.850 39.585 ;
        RECT 46.090 39.510 46.350 39.585 ;
        RECT 34.525 39.340 46.350 39.510 ;
        RECT 34.525 39.230 34.825 39.340 ;
        RECT 41.590 39.265 41.850 39.340 ;
        RECT 46.090 39.265 46.350 39.340 ;
        RECT 37.525 39.090 37.825 39.200 ;
        RECT 40.090 39.090 40.350 39.165 ;
        RECT 37.525 38.920 40.350 39.090 ;
        RECT 37.525 38.810 37.825 38.920 ;
        RECT 40.090 38.845 40.350 38.920 ;
        RECT 36.025 38.670 36.325 38.780 ;
        RECT 44.590 38.670 44.850 38.745 ;
        RECT 36.025 38.500 44.850 38.670 ;
        RECT 36.025 38.390 36.325 38.500 ;
        RECT 44.590 38.425 44.850 38.500 ;
        RECT 38.590 38.315 38.850 38.325 ;
        RECT 38.590 38.250 39.370 38.315 ;
        RECT 43.090 38.250 43.350 38.325 ;
        RECT 37.590 38.080 43.350 38.250 ;
        RECT 38.590 38.015 39.370 38.080 ;
        RECT 38.590 38.005 38.850 38.015 ;
        RECT 43.090 38.005 43.350 38.080 ;
        RECT 32.315 37.775 32.575 37.850 ;
        RECT 32.315 37.605 43.760 37.775 ;
        RECT 32.315 37.530 32.575 37.605 ;
        RECT 15.975 37.095 16.385 37.445 ;
        RECT 28.645 37.355 28.965 37.400 ;
        RECT 35.560 37.355 35.880 37.400 ;
        RECT 28.645 37.185 35.880 37.355 ;
        RECT 28.645 37.140 28.965 37.185 ;
        RECT 35.560 37.140 35.880 37.185 ;
        RECT 36.045 37.355 36.305 37.430 ;
        RECT 37.090 37.355 37.350 37.430 ;
        RECT 36.045 37.185 37.350 37.355 ;
        RECT 36.045 37.110 36.305 37.185 ;
        RECT 37.090 37.110 37.350 37.185 ;
        RECT 39.045 37.355 39.305 37.430 ;
        RECT 40.545 37.355 40.805 37.430 ;
        RECT 42.025 37.355 42.325 37.465 ;
        RECT 43.590 37.430 43.760 37.605 ;
        RECT 39.045 37.185 42.325 37.355 ;
        RECT 39.045 37.110 39.305 37.185 ;
        RECT 40.545 37.110 40.805 37.185 ;
        RECT 42.025 37.075 42.325 37.185 ;
        RECT 43.545 37.355 43.805 37.430 ;
        RECT 45.045 37.355 45.305 37.430 ;
        RECT 46.525 37.355 46.825 37.465 ;
        RECT 43.545 37.185 46.825 37.355 ;
        RECT 43.545 37.110 43.805 37.185 ;
        RECT 45.045 37.110 45.305 37.185 ;
        RECT 46.525 37.075 46.825 37.185 ;
        RECT 33.085 35.550 33.345 35.625 ;
        RECT 34.090 35.550 34.350 35.625 ;
        RECT 33.085 35.380 34.350 35.550 ;
        RECT 33.085 35.305 33.345 35.380 ;
        RECT 34.090 35.305 34.350 35.380 ;
        RECT 35.275 34.420 35.575 34.810 ;
        RECT 38.275 34.420 38.575 34.810 ;
        RECT 41.275 34.420 41.575 34.810 ;
        RECT 44.275 34.420 44.575 34.810 ;
        RECT 49.330 33.435 49.830 48.365 ;
        RECT 54.480 48.335 69.160 49.025 ;
        RECT 53.090 48.130 53.390 48.160 ;
        RECT 53.045 48.100 53.435 48.130 ;
        RECT 53.045 47.830 53.580 48.100 ;
        RECT 53.090 47.800 53.580 47.830 ;
        RECT 51.930 46.840 52.680 47.530 ;
        RECT 50.550 40.780 51.300 41.470 ;
        RECT 39.760 32.935 49.830 33.435 ;
        RECT 39.760 0.975 40.260 32.935 ;
        RECT 50.580 25.165 51.270 40.780 ;
        RECT 51.960 33.415 52.650 46.840 ;
        RECT 53.340 38.395 53.580 47.800 ;
        RECT 54.480 47.530 55.170 48.335 ;
        RECT 54.450 46.840 55.200 47.530 ;
        RECT 56.050 47.250 56.740 47.940 ;
        RECT 57.430 47.250 58.120 47.940 ;
        RECT 58.810 47.250 59.500 47.940 ;
        RECT 60.190 47.250 60.880 47.940 ;
        RECT 61.570 47.250 62.260 47.940 ;
        RECT 62.950 47.250 63.640 47.940 ;
        RECT 64.330 47.250 65.020 47.940 ;
        RECT 65.710 47.250 66.400 47.940 ;
        RECT 67.090 47.250 67.780 47.940 ;
        RECT 68.470 47.250 69.160 47.940 ;
        RECT 55.540 46.690 56.370 47.010 ;
        RECT 55.540 46.035 56.255 46.690 ;
        RECT 56.510 46.495 56.740 47.250 ;
        RECT 56.920 46.690 57.750 47.010 ;
        RECT 56.510 46.175 56.770 46.495 ;
        RECT 56.920 46.320 57.635 46.690 ;
        RECT 57.405 46.035 57.635 46.320 ;
        RECT 57.890 46.495 58.120 47.250 ;
        RECT 58.300 46.690 59.130 47.010 ;
        RECT 57.890 46.175 58.150 46.495 ;
        RECT 58.300 46.320 59.015 46.690 ;
        RECT 58.785 46.035 59.015 46.320 ;
        RECT 59.270 46.495 59.500 47.250 ;
        RECT 59.680 46.690 60.510 47.010 ;
        RECT 59.270 46.175 59.530 46.495 ;
        RECT 59.680 46.320 60.395 46.690 ;
        RECT 60.165 46.035 60.395 46.320 ;
        RECT 60.650 46.495 60.880 47.250 ;
        RECT 61.060 46.690 61.890 47.010 ;
        RECT 60.650 46.175 60.910 46.495 ;
        RECT 61.060 46.320 61.775 46.690 ;
        RECT 61.545 46.035 61.775 46.320 ;
        RECT 62.030 46.495 62.260 47.250 ;
        RECT 62.440 46.690 63.270 47.010 ;
        RECT 62.030 46.175 62.290 46.495 ;
        RECT 62.440 46.320 63.155 46.690 ;
        RECT 62.925 46.035 63.155 46.320 ;
        RECT 63.410 46.495 63.640 47.250 ;
        RECT 63.820 46.690 64.650 47.010 ;
        RECT 63.410 46.175 63.670 46.495 ;
        RECT 63.820 46.320 64.535 46.690 ;
        RECT 64.305 46.035 64.535 46.320 ;
        RECT 64.790 46.495 65.020 47.250 ;
        RECT 65.200 46.690 66.030 47.010 ;
        RECT 64.790 46.175 65.050 46.495 ;
        RECT 65.200 46.320 65.915 46.690 ;
        RECT 65.685 46.035 65.915 46.320 ;
        RECT 66.170 46.495 66.400 47.250 ;
        RECT 66.580 46.690 67.410 47.010 ;
        RECT 66.170 46.175 66.430 46.495 ;
        RECT 66.580 46.320 67.295 46.690 ;
        RECT 67.065 46.035 67.295 46.320 ;
        RECT 67.550 46.495 67.780 47.250 ;
        RECT 67.960 46.690 68.790 47.010 ;
        RECT 67.550 46.175 67.810 46.495 ;
        RECT 67.960 46.035 68.675 46.690 ;
        RECT 68.930 46.495 69.160 47.250 ;
        RECT 68.930 46.175 69.190 46.495 ;
        RECT 55.540 45.805 56.740 46.035 ;
        RECT 57.405 45.805 58.120 46.035 ;
        RECT 58.785 45.805 59.500 46.035 ;
        RECT 60.165 45.805 60.880 46.035 ;
        RECT 61.545 45.805 62.260 46.035 ;
        RECT 62.925 45.805 63.640 46.035 ;
        RECT 64.305 45.805 65.020 46.035 ;
        RECT 65.685 45.805 66.400 46.035 ;
        RECT 67.065 45.805 67.780 46.035 ;
        RECT 53.790 45.125 54.090 45.515 ;
        RECT 53.820 38.875 54.060 45.125 ;
        RECT 55.540 44.970 56.230 45.805 ;
        RECT 55.910 44.785 56.370 44.830 ;
        RECT 55.540 44.555 56.370 44.785 ;
        RECT 54.450 40.780 55.200 41.470 ;
        RECT 54.480 39.905 55.170 40.780 ;
        RECT 55.540 40.720 55.770 44.555 ;
        RECT 55.910 44.510 56.370 44.555 ;
        RECT 55.910 42.850 56.370 42.895 ;
        RECT 56.510 42.850 56.740 45.805 ;
        RECT 56.920 44.970 57.610 45.665 ;
        RECT 57.290 44.785 57.750 44.830 ;
        RECT 55.910 42.620 56.740 42.850 ;
        RECT 56.920 44.555 57.750 44.785 ;
        RECT 55.910 42.575 56.370 42.620 ;
        RECT 55.540 40.070 55.860 40.720 ;
        RECT 56.050 39.905 56.740 42.430 ;
        RECT 56.920 40.720 57.150 44.555 ;
        RECT 57.290 44.510 57.750 44.555 ;
        RECT 57.290 42.850 57.750 42.895 ;
        RECT 57.890 42.850 58.120 45.805 ;
        RECT 58.300 44.970 58.990 45.665 ;
        RECT 58.670 44.785 59.130 44.830 ;
        RECT 57.290 42.620 58.120 42.850 ;
        RECT 58.300 44.555 59.130 44.785 ;
        RECT 57.290 42.575 57.750 42.620 ;
        RECT 57.430 41.740 58.120 42.430 ;
        RECT 57.430 40.880 58.120 41.570 ;
        RECT 58.300 40.720 58.530 44.555 ;
        RECT 58.670 44.510 59.130 44.555 ;
        RECT 58.670 42.850 59.130 42.895 ;
        RECT 59.270 42.850 59.500 45.805 ;
        RECT 59.680 44.970 60.370 45.665 ;
        RECT 60.050 44.785 60.510 44.830 ;
        RECT 58.670 42.620 59.500 42.850 ;
        RECT 59.680 44.555 60.510 44.785 ;
        RECT 58.670 42.575 59.130 42.620 ;
        RECT 58.810 41.740 59.500 42.430 ;
        RECT 58.810 40.880 59.500 41.570 ;
        RECT 59.680 40.720 59.910 44.555 ;
        RECT 60.050 44.510 60.510 44.555 ;
        RECT 60.050 42.850 60.510 42.895 ;
        RECT 60.650 42.850 60.880 45.805 ;
        RECT 61.060 44.970 61.750 45.665 ;
        RECT 61.430 44.785 61.890 44.830 ;
        RECT 60.050 42.620 60.880 42.850 ;
        RECT 61.060 44.555 61.890 44.785 ;
        RECT 60.050 42.575 60.510 42.620 ;
        RECT 60.190 41.740 60.880 42.430 ;
        RECT 60.190 40.880 60.880 41.570 ;
        RECT 61.060 40.720 61.290 44.555 ;
        RECT 61.430 44.510 61.890 44.555 ;
        RECT 61.430 42.850 61.890 42.895 ;
        RECT 62.030 42.850 62.260 45.805 ;
        RECT 62.440 44.970 63.130 45.665 ;
        RECT 62.810 44.785 63.270 44.830 ;
        RECT 61.430 42.620 62.260 42.850 ;
        RECT 62.440 44.555 63.270 44.785 ;
        RECT 61.430 42.575 61.890 42.620 ;
        RECT 61.570 41.740 62.260 42.430 ;
        RECT 61.570 40.880 62.260 41.570 ;
        RECT 62.440 40.720 62.670 44.555 ;
        RECT 62.810 44.510 63.270 44.555 ;
        RECT 62.810 42.850 63.270 42.895 ;
        RECT 63.410 42.850 63.640 45.805 ;
        RECT 63.820 44.970 64.510 45.665 ;
        RECT 64.190 44.785 64.650 44.830 ;
        RECT 62.810 42.620 63.640 42.850 ;
        RECT 63.820 44.555 64.650 44.785 ;
        RECT 62.810 42.575 63.270 42.620 ;
        RECT 62.950 41.740 63.640 42.430 ;
        RECT 62.950 40.880 63.640 41.570 ;
        RECT 63.820 40.720 64.050 44.555 ;
        RECT 64.190 44.510 64.650 44.555 ;
        RECT 64.190 42.850 64.650 42.895 ;
        RECT 64.790 42.850 65.020 45.805 ;
        RECT 65.200 44.970 65.890 45.665 ;
        RECT 65.570 44.785 66.030 44.830 ;
        RECT 64.190 42.620 65.020 42.850 ;
        RECT 65.200 44.555 66.030 44.785 ;
        RECT 64.190 42.575 64.650 42.620 ;
        RECT 64.330 41.740 65.020 42.430 ;
        RECT 64.330 40.880 65.020 41.570 ;
        RECT 65.200 40.720 65.430 44.555 ;
        RECT 65.570 44.510 66.030 44.555 ;
        RECT 65.570 42.850 66.030 42.895 ;
        RECT 66.170 42.850 66.400 45.805 ;
        RECT 66.580 44.970 67.270 45.665 ;
        RECT 66.950 44.785 67.410 44.830 ;
        RECT 65.570 42.620 66.400 42.850 ;
        RECT 66.580 44.555 67.410 44.785 ;
        RECT 65.570 42.575 66.030 42.620 ;
        RECT 65.710 41.740 66.400 42.430 ;
        RECT 65.710 40.880 66.400 41.570 ;
        RECT 66.580 40.720 66.810 44.555 ;
        RECT 66.950 44.510 67.410 44.555 ;
        RECT 66.950 42.850 67.410 42.895 ;
        RECT 67.550 42.850 67.780 45.805 ;
        RECT 67.960 45.805 69.160 46.035 ;
        RECT 67.960 44.970 68.650 45.805 ;
        RECT 68.330 44.785 68.790 44.830 ;
        RECT 66.950 42.620 67.780 42.850 ;
        RECT 67.960 44.555 68.790 44.785 ;
        RECT 66.950 42.575 67.410 42.620 ;
        RECT 67.090 41.740 67.780 42.430 ;
        RECT 67.090 40.880 67.780 41.570 ;
        RECT 67.960 40.720 68.190 44.555 ;
        RECT 68.330 44.510 68.790 44.555 ;
        RECT 68.330 42.850 68.790 42.895 ;
        RECT 68.930 42.850 69.160 45.805 ;
        RECT 68.330 42.620 69.160 42.850 ;
        RECT 68.330 42.575 68.790 42.620 ;
        RECT 56.920 40.070 57.240 40.720 ;
        RECT 58.300 40.070 58.620 40.720 ;
        RECT 59.680 40.070 60.000 40.720 ;
        RECT 61.060 40.070 61.380 40.720 ;
        RECT 62.440 40.070 62.760 40.720 ;
        RECT 63.820 40.070 64.140 40.720 ;
        RECT 65.200 40.070 65.520 40.720 ;
        RECT 66.580 40.070 66.900 40.720 ;
        RECT 67.960 40.070 68.280 40.720 ;
        RECT 68.470 39.905 69.160 42.430 ;
        RECT 54.480 39.215 69.200 39.905 ;
        RECT 69.695 38.875 69.935 49.580 ;
        RECT 53.820 38.635 56.600 38.875 ;
        RECT 53.340 38.155 55.160 38.395 ;
        RECT 56.360 38.155 56.600 38.635 ;
        RECT 58.240 38.635 69.935 38.875 ;
        RECT 58.240 38.155 58.480 38.635 ;
        RECT 51.940 32.775 52.670 33.415 ;
        RECT 51.960 32.750 52.650 32.775 ;
        RECT 54.920 29.125 55.160 38.155 ;
        RECT 56.000 37.835 56.960 38.155 ;
        RECT 57.880 37.835 58.840 38.155 ;
        RECT 59.760 37.885 62.600 38.205 ;
        RECT 64.755 38.075 65.075 38.335 ;
        RECT 64.790 37.685 65.040 38.075 ;
        RECT 60.690 37.525 61.690 37.675 ;
        RECT 62.750 37.525 63.750 37.685 ;
        RECT 64.640 37.525 65.640 37.685 ;
        RECT 60.690 37.285 69.940 37.525 ;
        RECT 60.690 36.675 61.690 37.285 ;
        RECT 62.750 36.685 63.750 37.285 ;
        RECT 64.640 36.685 65.640 37.285 ;
        RECT 57.315 34.185 63.220 34.425 ;
        RECT 57.315 33.905 57.555 34.185 ;
        RECT 56.000 32.705 56.960 33.465 ;
        RECT 56.360 29.995 56.600 32.705 ;
        RECT 57.170 32.265 57.700 33.905 ;
        RECT 57.890 32.705 58.830 33.465 ;
        RECT 59.760 33.210 60.720 33.475 ;
        RECT 61.640 33.210 62.600 33.475 ;
        RECT 59.760 32.960 62.600 33.210 ;
        RECT 58.240 31.045 58.480 32.705 ;
        RECT 59.760 32.695 60.720 32.960 ;
        RECT 61.640 32.695 62.600 32.960 ;
        RECT 58.240 30.805 62.250 31.045 ;
        RECT 56.360 29.755 60.370 29.995 ;
        RECT 55.350 29.125 56.350 29.505 ;
        RECT 54.920 28.885 56.350 29.125 ;
        RECT 55.350 28.505 56.350 28.885 ;
        RECT 59.380 28.505 59.990 29.105 ;
        RECT 55.750 28.020 56.000 28.505 ;
        RECT 59.560 28.020 59.810 28.505 ;
        RECT 55.750 27.770 59.810 28.020 ;
        RECT 55.750 27.345 56.000 27.770 ;
        RECT 55.580 26.735 56.180 27.345 ;
        RECT 59.560 27.335 59.810 27.770 ;
        RECT 59.380 26.735 59.990 27.335 ;
        RECT 59.560 25.830 59.810 26.735 ;
        RECT 59.325 25.580 59.810 25.830 ;
        RECT 50.560 24.525 51.290 25.165 ;
        RECT 56.000 24.925 56.960 25.185 ;
        RECT 57.880 24.925 58.850 25.195 ;
        RECT 56.000 24.675 58.850 24.925 ;
        RECT 56.000 24.415 56.960 24.675 ;
        RECT 57.880 24.415 58.850 24.675 ;
        RECT 59.325 23.410 59.575 25.580 ;
        RECT 60.130 25.185 60.370 29.755 ;
        RECT 62.010 28.005 62.250 30.805 ;
        RECT 62.980 28.855 63.220 34.185 ;
        RECT 63.500 33.210 64.500 33.475 ;
        RECT 65.380 33.210 66.380 33.475 ;
        RECT 63.500 32.960 66.380 33.210 ;
        RECT 63.500 32.695 64.500 32.960 ;
        RECT 65.380 32.695 66.380 32.960 ;
        RECT 69.700 30.455 69.940 37.285 ;
        RECT 64.340 28.855 64.950 29.035 ;
        RECT 62.980 28.615 64.950 28.855 ;
        RECT 64.340 28.435 64.950 28.615 ;
        RECT 66.220 28.435 66.830 29.035 ;
        RECT 62.010 27.765 65.430 28.005 ;
        RECT 59.760 24.415 60.720 25.185 ;
        RECT 60.120 23.845 60.360 24.415 ;
        RECT 60.905 24.265 61.465 25.585 ;
        RECT 62.010 25.185 62.250 27.765 ;
        RECT 64.350 27.165 64.950 27.335 ;
        RECT 62.940 26.925 64.950 27.165 ;
        RECT 61.640 24.415 62.600 25.185 ;
        RECT 62.940 24.265 63.180 26.925 ;
        RECT 64.350 26.735 64.950 26.925 ;
        RECT 65.190 26.355 65.430 27.765 ;
        RECT 66.405 27.335 66.655 28.435 ;
        RECT 69.640 28.235 69.990 30.455 ;
        RECT 74.350 29.910 74.700 120.295 ;
        RECT 112.700 120.250 113.050 177.705 ;
        RECT 113.310 176.775 113.610 176.840 ;
        RECT 113.300 176.515 113.620 176.775 ;
        RECT 113.310 176.450 113.610 176.515 ;
        RECT 114.200 118.750 114.550 177.705 ;
        RECT 114.810 176.775 115.110 176.840 ;
        RECT 114.800 176.515 115.120 176.775 ;
        RECT 114.810 176.450 115.110 176.515 ;
        RECT 115.700 117.250 116.050 177.705 ;
        RECT 116.310 176.775 116.610 176.840 ;
        RECT 116.300 176.515 116.620 176.775 ;
        RECT 116.310 176.450 116.610 176.515 ;
        RECT 117.200 115.750 117.550 177.705 ;
        RECT 117.810 176.775 118.110 176.840 ;
        RECT 117.800 176.515 118.120 176.775 ;
        RECT 117.810 176.450 118.110 176.515 ;
        RECT 118.700 114.250 119.050 177.705 ;
        RECT 119.435 176.790 119.735 176.840 ;
        RECT 119.410 176.500 119.760 176.790 ;
        RECT 119.435 176.450 119.735 176.500 ;
        RECT 89.900 104.700 93.820 104.980 ;
        RECT 87.380 104.420 96.060 104.700 ;
        RECT 85.420 104.140 97.180 104.420 ;
        RECT 84.300 103.860 98.300 104.140 ;
        RECT 83.460 103.580 99.140 103.860 ;
        RECT 82.900 103.300 99.700 103.580 ;
        RECT 82.340 103.020 100.540 103.300 ;
        RECT 81.780 102.740 101.100 103.020 ;
        RECT 81.500 102.460 101.380 102.740 ;
        RECT 80.940 102.180 101.940 102.460 ;
        RECT 80.660 101.900 102.500 102.180 ;
        RECT 80.380 101.620 102.780 101.900 ;
        RECT 80.100 101.340 89.060 101.620 ;
        RECT 94.380 101.340 103.060 101.620 ;
        RECT 80.100 101.060 87.380 101.340 ;
        RECT 96.340 101.060 103.340 101.340 ;
        RECT 79.820 100.780 85.980 101.060 ;
        RECT 97.180 100.780 103.620 101.060 ;
        RECT 79.540 100.500 85.420 100.780 ;
        RECT 98.020 100.500 103.620 100.780 ;
        RECT 79.540 100.220 84.860 100.500 ;
        RECT 98.300 100.220 103.900 100.500 ;
        RECT 79.540 99.940 84.580 100.220 ;
        RECT 98.580 99.940 103.900 100.220 ;
        RECT 79.260 99.660 84.580 99.940 ;
        RECT 98.860 99.660 103.900 99.940 ;
        RECT 79.260 97.420 84.300 99.660 ;
        RECT 86.540 99.380 88.220 99.660 ;
        RECT 94.940 99.380 96.620 99.660 ;
        RECT 85.980 99.100 88.500 99.380 ;
        RECT 94.660 99.100 97.180 99.380 ;
        RECT 85.980 98.820 88.780 99.100 ;
        RECT 94.660 98.820 97.460 99.100 ;
        RECT 85.700 98.540 88.780 98.820 ;
        RECT 85.700 97.980 89.060 98.540 ;
        RECT 94.380 98.260 97.460 98.820 ;
        RECT 89.900 97.980 93.260 98.260 ;
        RECT 94.100 97.980 97.460 98.260 ;
        RECT 85.980 97.420 97.180 97.980 ;
        RECT 79.540 97.140 84.300 97.420 ;
        RECT 79.540 96.580 84.020 97.140 ;
        RECT 86.260 96.860 97.180 97.420 ;
        RECT 98.860 97.420 104.180 99.660 ;
        RECT 98.860 97.140 103.900 97.420 ;
        RECT 99.140 96.860 103.900 97.140 ;
        RECT 79.820 96.300 83.460 96.580 ;
        RECT 85.980 96.300 97.460 96.860 ;
        RECT 99.420 96.580 103.620 96.860 ;
        RECT 99.700 96.300 103.340 96.580 ;
        RECT 80.100 96.020 82.900 96.300 ;
        RECT 80.660 95.740 82.340 96.020 ;
        RECT 85.700 95.740 97.740 96.300 ;
        RECT 100.540 96.020 102.780 96.300 ;
        RECT 85.420 95.460 91.020 95.740 ;
        RECT 92.700 95.460 98.020 95.740 ;
        RECT 85.140 95.180 90.180 95.460 ;
        RECT 93.540 95.180 98.300 95.460 ;
        RECT 85.140 94.900 89.620 95.180 ;
        RECT 94.100 94.900 98.300 95.180 ;
        RECT 84.860 94.620 89.060 94.900 ;
        RECT 94.660 94.620 98.580 94.900 ;
        RECT 84.580 94.340 88.780 94.620 ;
        RECT 94.940 94.340 98.580 94.620 ;
        RECT 84.580 94.060 88.500 94.340 ;
        RECT 95.220 94.060 98.860 94.340 ;
        RECT 84.300 93.780 88.220 94.060 ;
        RECT 84.020 93.500 88.220 93.780 ;
        RECT 90.740 93.500 92.980 93.780 ;
        RECT 95.500 93.500 99.140 94.060 ;
        RECT 84.020 93.220 87.940 93.500 ;
        RECT 90.180 93.220 93.260 93.500 ;
        RECT 83.740 92.660 87.660 93.220 ;
        RECT 89.900 92.940 93.540 93.220 ;
        RECT 95.780 92.940 99.420 93.500 ;
        RECT 83.460 92.380 87.660 92.660 ;
        RECT 89.620 92.380 93.820 92.940 ;
        RECT 96.060 92.380 99.700 92.940 ;
        RECT 83.460 92.100 87.380 92.380 ;
        RECT 83.180 91.820 87.380 92.100 ;
        RECT 82.900 91.260 87.380 91.820 ;
        RECT 82.620 90.700 87.380 91.260 ;
        RECT 89.340 90.980 94.100 92.380 ;
        RECT 96.060 91.540 99.980 92.380 ;
        RECT 96.060 90.980 100.260 91.540 ;
        RECT 82.340 90.140 87.660 90.700 ;
        RECT 89.620 90.420 93.820 90.980 ;
        RECT 96.060 90.700 100.540 90.980 ;
        RECT 95.780 90.420 100.540 90.700 ;
        RECT 89.900 90.140 93.540 90.420 ;
        RECT 95.780 90.140 100.820 90.420 ;
        RECT 82.060 89.860 87.660 90.140 ;
        RECT 90.180 89.860 93.260 90.140 ;
        RECT 82.060 89.300 87.940 89.860 ;
        RECT 90.740 89.580 92.700 89.860 ;
        RECT 95.500 89.580 100.820 90.140 ;
        RECT 81.780 89.020 88.220 89.300 ;
        RECT 95.220 89.020 101.100 89.580 ;
        RECT 81.780 88.740 88.500 89.020 ;
        RECT 94.940 88.740 101.380 89.020 ;
        RECT 81.500 88.460 88.780 88.740 ;
        RECT 94.660 88.460 101.380 88.740 ;
        RECT 81.500 88.180 89.060 88.460 ;
        RECT 94.100 88.180 101.380 88.460 ;
        RECT 81.500 87.900 89.620 88.180 ;
        RECT 93.820 87.900 101.380 88.180 ;
        RECT 81.220 87.620 90.180 87.900 ;
        RECT 92.980 87.620 101.660 87.900 ;
        RECT 81.220 85.100 101.660 87.620 ;
        RECT 81.780 84.820 101.100 85.100 ;
        RECT 108.385 41.385 136.870 41.885 ;
        RECT 102.225 38.950 102.575 41.110 ;
        RECT 108.385 40.530 108.885 41.385 ;
        RECT 108.125 39.530 109.125 40.530 ;
        RECT 114.735 39.560 115.795 40.500 ;
        RECT 102.280 38.755 102.520 38.950 ;
        RECT 115.140 38.755 115.385 39.560 ;
        RECT 121.315 38.950 121.665 41.110 ;
        RECT 121.365 38.755 121.605 38.950 ;
        RECT 102.280 38.515 113.975 38.755 ;
        RECT 107.140 38.075 107.460 38.335 ;
        RECT 107.175 37.685 107.425 38.075 ;
        RECT 109.615 37.885 112.455 38.205 ;
        RECT 113.735 38.155 113.975 38.515 ;
        RECT 115.140 38.510 115.860 38.755 ;
        RECT 116.625 38.515 121.605 38.755 ;
        RECT 115.615 38.155 115.855 38.510 ;
        RECT 113.375 37.835 114.335 38.155 ;
        RECT 115.255 37.835 116.215 38.155 ;
        RECT 106.575 37.525 107.575 37.685 ;
        RECT 108.465 37.525 109.465 37.685 ;
        RECT 110.525 37.525 111.525 37.675 ;
        RECT 102.275 37.285 111.525 37.525 ;
        RECT 86.770 31.360 87.460 32.140 ;
        RECT 86.770 30.320 87.460 31.010 ;
        RECT 102.275 30.455 102.515 37.285 ;
        RECT 106.575 36.685 107.575 37.285 ;
        RECT 108.465 36.685 109.465 37.285 ;
        RECT 110.525 36.675 111.525 37.285 ;
        RECT 108.995 34.185 114.900 34.425 ;
        RECT 105.835 33.210 106.835 33.475 ;
        RECT 107.715 33.210 108.715 33.475 ;
        RECT 105.835 32.960 108.715 33.210 ;
        RECT 105.835 32.695 106.835 32.960 ;
        RECT 107.715 32.695 108.715 32.960 ;
        RECT 86.260 29.910 87.090 30.080 ;
        RECT 74.350 29.905 84.450 29.910 ;
        RECT 85.455 29.905 87.090 29.910 ;
        RECT 74.350 29.760 87.090 29.905 ;
        RECT 74.350 29.560 86.975 29.760 ;
        RECT 86.260 29.390 86.975 29.560 ;
        RECT 86.745 29.105 86.975 29.390 ;
        RECT 87.230 29.565 87.460 30.320 ;
        RECT 87.230 29.245 87.490 29.565 ;
        RECT 86.745 28.875 87.460 29.105 ;
        RECT 86.260 28.635 86.950 28.735 ;
        RECT 69.690 27.915 69.940 28.235 ;
        RECT 84.595 28.135 86.950 28.635 ;
        RECT 66.230 26.735 66.830 27.335 ;
        RECT 68.990 26.915 69.990 27.915 ;
        RECT 68.990 26.375 69.990 26.625 ;
        RECT 84.595 26.375 85.095 28.135 ;
        RECT 86.260 28.040 86.950 28.135 ;
        RECT 86.630 27.855 87.090 27.900 ;
        RECT 68.990 26.355 85.095 26.375 ;
        RECT 65.190 26.115 85.095 26.355 ;
        RECT 68.990 25.875 85.095 26.115 ;
        RECT 86.260 27.625 87.090 27.855 ;
        RECT 68.990 25.625 69.990 25.875 ;
        RECT 63.500 24.925 64.500 25.185 ;
        RECT 65.380 24.925 66.380 25.185 ;
        RECT 67.260 24.925 68.260 25.185 ;
        RECT 63.500 24.675 68.260 24.925 ;
        RECT 68.990 24.805 69.990 25.345 ;
        RECT 63.500 24.415 64.500 24.675 ;
        RECT 65.380 24.415 66.380 24.675 ;
        RECT 67.260 24.415 68.260 24.675 ;
        RECT 68.550 24.565 69.990 24.805 ;
        RECT 60.905 24.025 63.180 24.265 ;
        RECT 68.550 23.845 68.790 24.565 ;
        RECT 68.990 24.345 69.990 24.565 ;
        RECT 60.120 23.605 68.790 23.845 ;
        RECT 68.990 23.795 69.990 24.045 ;
        RECT 68.990 23.410 71.305 23.795 ;
        RECT 59.325 23.295 71.305 23.410 ;
        RECT 59.325 23.160 69.990 23.295 ;
        RECT 68.990 23.045 69.990 23.160 ;
        RECT 56.770 22.705 58.090 23.035 ;
        RECT 62.810 22.705 64.130 23.015 ;
        RECT 64.690 22.705 66.010 23.015 ;
        RECT 66.570 22.705 67.890 23.005 ;
        RECT 68.990 22.735 69.990 22.775 ;
        RECT 68.700 22.705 69.990 22.735 ;
        RECT 56.770 22.465 69.990 22.705 ;
        RECT 56.770 22.275 58.090 22.465 ;
        RECT 62.810 22.255 64.130 22.465 ;
        RECT 64.690 22.255 66.010 22.465 ;
        RECT 66.570 22.245 67.890 22.465 ;
        RECT 55.990 22.105 56.980 22.135 ;
        RECT 57.860 22.105 58.840 22.135 ;
        RECT 55.990 21.855 58.840 22.105 ;
        RECT 55.990 21.815 56.980 21.855 ;
        RECT 57.860 21.815 58.840 21.855 ;
        RECT 63.500 22.060 64.500 22.095 ;
        RECT 65.380 22.060 66.380 22.095 ;
        RECT 67.260 22.060 68.260 22.095 ;
        RECT 63.500 21.810 68.260 22.060 ;
        RECT 63.500 21.775 64.500 21.810 ;
        RECT 65.380 21.775 66.380 21.810 ;
        RECT 67.260 21.775 68.260 21.810 ;
        RECT 68.990 21.775 69.990 22.465 ;
        RECT 70.805 18.585 71.305 23.295 ;
        RECT 59.085 18.085 71.305 18.585 ;
        RECT 59.085 0.975 59.585 18.085 ;
        RECT 78.395 0.975 78.895 25.875 ;
        RECT 86.260 23.790 86.490 27.625 ;
        RECT 86.630 27.580 87.090 27.625 ;
        RECT 86.630 25.920 87.090 25.965 ;
        RECT 87.230 25.920 87.460 28.875 ;
        RECT 102.225 28.235 102.575 30.455 ;
        RECT 105.385 28.435 105.995 29.035 ;
        RECT 107.265 28.855 107.875 29.035 ;
        RECT 108.995 28.855 109.235 34.185 ;
        RECT 114.660 33.905 114.900 34.185 ;
        RECT 109.615 33.210 110.575 33.475 ;
        RECT 111.495 33.210 112.455 33.475 ;
        RECT 109.615 32.960 112.455 33.210 ;
        RECT 109.615 32.695 110.575 32.960 ;
        RECT 111.495 32.695 112.455 32.960 ;
        RECT 113.385 32.705 114.325 33.465 ;
        RECT 113.735 31.045 113.975 32.705 ;
        RECT 114.515 32.265 115.045 33.905 ;
        RECT 115.255 32.705 116.215 33.465 ;
        RECT 107.265 28.615 109.235 28.855 ;
        RECT 109.965 30.805 113.975 31.045 ;
        RECT 107.265 28.435 107.875 28.615 ;
        RECT 102.275 27.915 102.525 28.235 ;
        RECT 102.225 26.915 103.225 27.915 ;
        RECT 105.560 27.335 105.810 28.435 ;
        RECT 109.965 28.005 110.205 30.805 ;
        RECT 115.615 29.995 115.855 32.705 ;
        RECT 106.785 27.765 110.205 28.005 ;
        RECT 105.385 26.735 105.985 27.335 ;
        RECT 102.225 26.375 103.225 26.625 ;
        RECT 86.630 25.690 87.460 25.920 ;
        RECT 88.555 26.355 103.225 26.375 ;
        RECT 106.785 26.355 107.025 27.765 ;
        RECT 107.265 27.165 107.865 27.335 ;
        RECT 107.265 26.925 109.275 27.165 ;
        RECT 107.265 26.735 107.865 26.925 ;
        RECT 88.555 26.115 107.025 26.355 ;
        RECT 88.555 25.875 103.225 26.115 ;
        RECT 86.630 25.645 87.090 25.690 ;
        RECT 86.770 25.405 87.460 25.500 ;
        RECT 88.555 25.405 89.055 25.875 ;
        RECT 86.770 24.905 89.055 25.405 ;
        RECT 86.770 24.810 87.460 24.905 ;
        RECT 86.770 23.950 87.460 24.640 ;
        RECT 86.260 23.140 86.580 23.790 ;
        RECT 86.770 22.240 87.460 23.020 ;
        RECT 97.740 0.975 98.240 25.875 ;
        RECT 102.225 25.625 103.225 25.875 ;
        RECT 102.225 24.805 103.225 25.345 ;
        RECT 103.955 24.925 104.955 25.185 ;
        RECT 105.835 24.925 106.835 25.185 ;
        RECT 107.715 24.925 108.715 25.185 ;
        RECT 102.225 24.565 103.665 24.805 ;
        RECT 102.225 24.345 103.225 24.565 ;
        RECT 102.225 23.795 103.225 24.045 ;
        RECT 101.225 23.410 103.225 23.795 ;
        RECT 103.425 23.845 103.665 24.565 ;
        RECT 103.955 24.675 108.715 24.925 ;
        RECT 103.955 24.415 104.955 24.675 ;
        RECT 105.835 24.415 106.835 24.675 ;
        RECT 107.715 24.415 108.715 24.675 ;
        RECT 109.035 24.265 109.275 26.925 ;
        RECT 109.965 25.185 110.205 27.765 ;
        RECT 111.845 29.755 115.855 29.995 ;
        RECT 109.615 24.415 110.575 25.185 ;
        RECT 110.750 24.265 111.310 25.585 ;
        RECT 111.845 25.185 112.085 29.755 ;
        RECT 116.625 29.505 116.865 38.515 ;
        RECT 112.225 28.505 112.835 29.105 ;
        RECT 115.865 28.505 116.865 29.505 ;
        RECT 112.405 28.020 112.655 28.505 ;
        RECT 116.215 28.020 116.465 28.505 ;
        RECT 112.405 27.770 116.465 28.020 ;
        RECT 112.405 27.335 112.655 27.770 ;
        RECT 116.215 27.345 116.465 27.770 ;
        RECT 112.225 26.735 112.835 27.335 ;
        RECT 116.035 26.735 116.635 27.345 ;
        RECT 112.405 25.830 112.655 26.735 ;
        RECT 112.405 25.580 112.890 25.830 ;
        RECT 111.495 24.415 112.455 25.185 ;
        RECT 109.035 24.025 111.310 24.265 ;
        RECT 111.855 23.845 112.095 24.415 ;
        RECT 103.425 23.605 112.095 23.845 ;
        RECT 112.640 23.410 112.890 25.580 ;
        RECT 113.365 24.925 114.335 25.195 ;
        RECT 115.255 24.925 116.215 25.185 ;
        RECT 113.365 24.675 116.215 24.925 ;
        RECT 113.365 24.415 114.335 24.675 ;
        RECT 115.255 24.415 116.215 24.675 ;
        RECT 101.225 23.295 112.890 23.410 ;
        RECT 101.225 18.615 101.725 23.295 ;
        RECT 102.225 23.160 112.890 23.295 ;
        RECT 102.225 23.045 103.225 23.160 ;
        RECT 102.225 22.735 103.225 22.775 ;
        RECT 102.225 22.705 103.515 22.735 ;
        RECT 104.325 22.705 105.645 23.005 ;
        RECT 106.205 22.705 107.525 23.015 ;
        RECT 108.085 22.705 109.405 23.015 ;
        RECT 114.125 22.705 115.445 23.035 ;
        RECT 102.225 22.465 115.445 22.705 ;
        RECT 102.225 21.775 103.225 22.465 ;
        RECT 104.325 22.245 105.645 22.465 ;
        RECT 106.205 22.255 107.525 22.465 ;
        RECT 108.085 22.255 109.405 22.465 ;
        RECT 114.125 22.275 115.445 22.465 ;
        RECT 113.375 22.105 114.355 22.135 ;
        RECT 115.235 22.105 116.225 22.135 ;
        RECT 103.955 22.060 104.955 22.095 ;
        RECT 105.835 22.060 106.835 22.095 ;
        RECT 107.715 22.060 108.715 22.095 ;
        RECT 103.955 21.810 108.715 22.060 ;
        RECT 113.375 21.855 116.225 22.105 ;
        RECT 113.375 21.815 114.355 21.855 ;
        RECT 115.235 21.815 116.225 21.855 ;
        RECT 103.955 21.775 104.955 21.810 ;
        RECT 105.835 21.775 106.835 21.810 ;
        RECT 107.715 21.775 108.715 21.810 ;
        RECT 101.225 18.115 117.555 18.615 ;
        RECT 117.055 0.975 117.555 18.115 ;
        RECT 136.370 0.975 136.870 41.385 ;
        RECT 39.550 0.125 40.490 0.975 ;
        RECT 58.870 0.125 59.810 0.975 ;
        RECT 78.190 0.125 79.130 0.975 ;
        RECT 97.510 0.125 98.450 0.975 ;
        RECT 116.830 0.125 117.770 0.975 ;
        RECT 136.150 0.125 137.090 0.975 ;
      LAYER met3 ;
        RECT 15.005 225.080 15.355 225.085 ;
        RECT 17.765 225.080 18.115 225.085 ;
        RECT 20.525 225.080 20.875 225.085 ;
        RECT 23.285 225.080 23.635 225.085 ;
        RECT 26.045 225.080 26.395 225.085 ;
        RECT 28.805 225.080 29.155 225.085 ;
        RECT 31.565 225.080 31.915 225.085 ;
        RECT 34.325 225.080 34.675 225.085 ;
        RECT 37.085 225.080 37.435 225.085 ;
        RECT 39.845 225.080 40.195 225.085 ;
        RECT 42.605 225.080 42.955 225.085 ;
        RECT 45.365 225.080 45.715 225.085 ;
        RECT 48.125 225.080 48.475 225.085 ;
        RECT 50.885 225.080 51.235 225.085 ;
        RECT 53.645 225.080 53.995 225.085 ;
        RECT 56.405 225.080 56.755 225.085 ;
        RECT 59.165 225.080 59.515 225.085 ;
        RECT 61.925 225.080 62.275 225.085 ;
        RECT 64.685 225.080 65.035 225.085 ;
        RECT 67.445 225.080 67.795 225.085 ;
        RECT 70.205 225.080 70.555 225.085 ;
        RECT 72.965 225.080 73.315 225.085 ;
        RECT 75.725 225.080 76.075 225.085 ;
        RECT 78.485 225.080 78.835 225.085 ;
        RECT 103.325 225.080 103.675 225.085 ;
        RECT 106.085 225.080 106.435 225.085 ;
        RECT 108.845 225.080 109.195 225.085 ;
        RECT 111.605 225.080 111.955 225.085 ;
        RECT 114.365 225.080 114.715 225.085 ;
        RECT 117.125 225.080 117.475 225.085 ;
        RECT 119.885 225.080 120.235 225.085 ;
        RECT 122.645 225.080 122.995 225.085 ;
        RECT 14.980 224.740 15.380 225.080 ;
        RECT 17.740 224.740 18.140 225.080 ;
        RECT 20.500 224.740 20.900 225.080 ;
        RECT 23.260 224.740 23.660 225.080 ;
        RECT 26.020 224.740 26.420 225.080 ;
        RECT 28.780 224.740 29.180 225.080 ;
        RECT 31.540 224.740 31.940 225.080 ;
        RECT 34.300 224.740 34.700 225.080 ;
        RECT 37.060 224.740 37.460 225.080 ;
        RECT 39.820 224.740 40.220 225.080 ;
        RECT 42.580 224.740 42.980 225.080 ;
        RECT 45.340 224.740 45.740 225.080 ;
        RECT 48.100 224.740 48.500 225.080 ;
        RECT 50.860 224.740 51.260 225.080 ;
        RECT 53.620 224.740 54.020 225.080 ;
        RECT 56.380 224.740 56.780 225.080 ;
        RECT 59.140 224.740 59.540 225.080 ;
        RECT 61.900 224.740 62.300 225.080 ;
        RECT 64.660 224.740 65.060 225.080 ;
        RECT 67.420 224.740 67.820 225.080 ;
        RECT 70.180 224.740 70.580 225.080 ;
        RECT 72.940 224.740 73.340 225.080 ;
        RECT 75.700 224.740 76.100 225.080 ;
        RECT 78.460 224.740 78.860 225.080 ;
        RECT 103.300 224.740 103.700 225.080 ;
        RECT 106.060 224.740 106.460 225.080 ;
        RECT 108.820 224.740 109.220 225.080 ;
        RECT 111.580 224.740 111.980 225.080 ;
        RECT 114.340 224.740 114.740 225.080 ;
        RECT 117.100 224.740 117.500 225.080 ;
        RECT 119.860 224.740 120.260 225.080 ;
        RECT 122.620 224.740 123.020 225.080 ;
        RECT 15.005 223.035 15.355 224.740 ;
        RECT 17.765 223.035 18.115 224.740 ;
        RECT 20.525 223.035 20.875 224.740 ;
        RECT 23.285 223.035 23.635 224.740 ;
        RECT 26.045 223.035 26.395 224.740 ;
        RECT 28.805 223.035 29.155 224.740 ;
        RECT 31.565 223.035 31.915 224.740 ;
        RECT 34.325 223.035 34.675 224.740 ;
        RECT 37.085 223.035 37.435 224.740 ;
        RECT 39.845 223.035 40.195 224.740 ;
        RECT 42.605 223.035 42.955 224.740 ;
        RECT 45.365 223.035 45.715 224.740 ;
        RECT 48.125 223.035 48.475 224.740 ;
        RECT 50.885 223.035 51.235 224.740 ;
        RECT 53.645 223.035 53.995 224.740 ;
        RECT 56.405 223.035 56.755 224.740 ;
        RECT 59.165 223.035 59.515 224.740 ;
        RECT 61.925 223.035 62.275 224.740 ;
        RECT 64.685 223.035 65.035 224.740 ;
        RECT 67.445 223.035 67.795 224.740 ;
        RECT 70.205 223.035 70.555 224.740 ;
        RECT 72.965 223.035 73.315 224.740 ;
        RECT 75.725 223.035 76.075 224.740 ;
        RECT 78.485 223.035 78.835 224.740 ;
        RECT 103.325 223.035 103.675 224.740 ;
        RECT 106.085 223.035 106.435 224.740 ;
        RECT 108.845 223.035 109.195 224.740 ;
        RECT 111.605 223.035 111.955 224.740 ;
        RECT 114.365 223.035 114.715 224.740 ;
        RECT 117.125 223.035 117.475 224.740 ;
        RECT 119.885 223.035 120.235 224.740 ;
        RECT 122.645 223.035 122.995 224.740 ;
        RECT 39.000 208.185 41.000 208.190 ;
        RECT 44.000 208.185 46.000 208.190 ;
        RECT 49.000 208.185 51.000 208.190 ;
        RECT 65.000 208.185 67.000 208.190 ;
        RECT 70.000 208.185 72.000 208.190 ;
        RECT 75.000 208.185 77.000 208.190 ;
        RECT 38.555 207.785 51.735 208.185 ;
        RECT 64.555 207.785 77.735 208.185 ;
        RECT 39.000 207.780 41.000 207.785 ;
        RECT 44.000 207.780 46.000 207.785 ;
        RECT 49.000 207.780 51.000 207.785 ;
        RECT 65.000 207.780 67.000 207.785 ;
        RECT 70.000 207.780 72.000 207.785 ;
        RECT 75.000 207.780 77.000 207.785 ;
        RECT 21.000 206.735 23.000 206.765 ;
        RECT 13.295 206.385 24.145 206.735 ;
        RECT 107.000 206.655 109.000 206.685 ;
        RECT 112.000 206.655 114.000 206.685 ;
        RECT 117.000 206.655 119.000 206.685 ;
        RECT 21.000 206.355 23.000 206.385 ;
        RECT 106.730 206.305 119.610 206.655 ;
        RECT 107.000 206.275 109.000 206.305 ;
        RECT 112.000 206.275 114.000 206.305 ;
        RECT 117.000 206.275 119.000 206.305 ;
        RECT 39.000 202.525 41.000 202.530 ;
        RECT 44.000 202.525 46.000 202.530 ;
        RECT 49.000 202.525 51.000 202.530 ;
        RECT 65.000 202.525 67.000 202.530 ;
        RECT 70.000 202.525 72.000 202.530 ;
        RECT 75.000 202.525 77.000 202.530 ;
        RECT 38.695 202.125 51.635 202.525 ;
        RECT 64.695 202.125 77.635 202.525 ;
        RECT 39.000 202.120 41.000 202.125 ;
        RECT 44.000 202.120 46.000 202.125 ;
        RECT 49.000 202.120 51.000 202.125 ;
        RECT 65.000 202.120 67.000 202.125 ;
        RECT 70.000 202.120 72.000 202.125 ;
        RECT 75.000 202.120 77.000 202.125 ;
        RECT 39.000 201.475 41.000 201.480 ;
        RECT 44.000 201.475 46.000 201.480 ;
        RECT 49.000 201.475 51.000 201.480 ;
        RECT 65.000 201.475 67.000 201.480 ;
        RECT 70.000 201.475 72.000 201.480 ;
        RECT 75.000 201.475 77.000 201.480 ;
        RECT 16.000 201.075 18.010 201.100 ;
        RECT 38.555 201.075 51.735 201.475 ;
        RECT 64.555 201.075 77.735 201.475 ;
        RECT 13.290 200.725 24.140 201.075 ;
        RECT 39.000 201.070 41.000 201.075 ;
        RECT 44.000 201.070 46.000 201.075 ;
        RECT 49.000 201.070 51.000 201.075 ;
        RECT 65.000 201.070 67.000 201.075 ;
        RECT 70.000 201.070 72.000 201.075 ;
        RECT 75.000 201.070 77.000 201.075 ;
        RECT 107.000 200.995 109.000 201.025 ;
        RECT 112.000 200.995 114.000 201.025 ;
        RECT 117.000 200.995 119.000 201.025 ;
        RECT 16.000 200.690 18.010 200.725 ;
        RECT 106.630 200.645 119.760 200.995 ;
        RECT 107.000 200.615 109.000 200.645 ;
        RECT 112.000 200.615 114.000 200.645 ;
        RECT 117.000 200.615 119.000 200.645 ;
        RECT 39.000 195.815 41.000 195.820 ;
        RECT 44.000 195.815 46.000 195.820 ;
        RECT 49.000 195.815 51.000 195.820 ;
        RECT 65.000 195.815 67.000 195.820 ;
        RECT 70.000 195.815 72.000 195.820 ;
        RECT 75.000 195.815 77.000 195.820 ;
        RECT 38.695 195.415 51.635 195.815 ;
        RECT 64.695 195.415 77.635 195.815 ;
        RECT 39.000 195.410 41.000 195.415 ;
        RECT 44.000 195.410 46.000 195.415 ;
        RECT 49.000 195.410 51.000 195.415 ;
        RECT 65.000 195.410 67.000 195.415 ;
        RECT 70.000 195.410 72.000 195.415 ;
        RECT 75.000 195.410 77.000 195.415 ;
        RECT 107.000 189.190 109.000 189.220 ;
        RECT 112.000 189.190 114.000 189.220 ;
        RECT 117.000 189.190 119.000 189.220 ;
        RECT 106.730 188.840 119.610 189.190 ;
        RECT 107.000 188.810 109.000 188.840 ;
        RECT 112.000 188.810 114.000 188.840 ;
        RECT 117.000 188.810 119.000 188.840 ;
        RECT 39.000 184.010 41.000 184.015 ;
        RECT 44.000 184.010 46.000 184.015 ;
        RECT 49.000 184.010 51.000 184.015 ;
        RECT 65.000 184.010 67.000 184.015 ;
        RECT 70.000 184.010 72.000 184.015 ;
        RECT 75.000 184.010 77.000 184.015 ;
        RECT 38.555 183.610 51.735 184.010 ;
        RECT 64.555 183.610 77.735 184.010 ;
        RECT 39.000 183.605 41.000 183.610 ;
        RECT 44.000 183.605 46.000 183.610 ;
        RECT 49.000 183.605 51.000 183.610 ;
        RECT 65.000 183.605 67.000 183.610 ;
        RECT 70.000 183.605 72.000 183.610 ;
        RECT 75.000 183.605 77.000 183.610 ;
        RECT 107.000 183.555 109.000 183.560 ;
        RECT 112.000 183.555 114.000 183.560 ;
        RECT 117.000 183.555 119.000 183.560 ;
        RECT 106.605 183.155 119.785 183.555 ;
        RECT 107.000 183.150 109.000 183.155 ;
        RECT 112.000 183.150 114.000 183.155 ;
        RECT 117.000 183.150 119.000 183.155 ;
        RECT 107.000 182.505 109.000 182.510 ;
        RECT 112.000 182.505 114.000 182.510 ;
        RECT 117.000 182.505 119.000 182.510 ;
        RECT 106.705 182.105 119.640 182.505 ;
        RECT 107.000 182.100 109.000 182.105 ;
        RECT 112.000 182.100 114.000 182.105 ;
        RECT 117.000 182.100 119.000 182.105 ;
        RECT 39.000 178.350 41.000 178.355 ;
        RECT 44.000 178.350 46.000 178.355 ;
        RECT 49.000 178.350 51.000 178.355 ;
        RECT 65.000 178.350 67.000 178.355 ;
        RECT 70.000 178.350 72.000 178.355 ;
        RECT 75.000 178.350 77.000 178.355 ;
        RECT 38.695 177.950 51.635 178.350 ;
        RECT 64.695 177.950 77.635 178.350 ;
        RECT 39.000 177.945 41.000 177.950 ;
        RECT 44.000 177.945 46.000 177.950 ;
        RECT 49.000 177.945 51.000 177.950 ;
        RECT 65.000 177.945 67.000 177.950 ;
        RECT 70.000 177.945 72.000 177.950 ;
        RECT 75.000 177.945 77.000 177.950 ;
        RECT 107.000 176.845 109.000 176.850 ;
        RECT 112.000 176.845 114.000 176.850 ;
        RECT 117.000 176.845 119.000 176.850 ;
        RECT 106.605 176.445 119.785 176.845 ;
        RECT 107.000 176.440 109.000 176.445 ;
        RECT 112.000 176.440 114.000 176.445 ;
        RECT 117.000 176.440 119.000 176.445 ;
        RECT 29.735 146.770 30.085 146.795 ;
        RECT 36.445 146.770 36.795 146.795 ;
        RECT 43.155 146.770 43.505 146.795 ;
        RECT 49.865 146.770 50.215 146.795 ;
        RECT 56.575 146.770 56.925 146.795 ;
        RECT 63.285 146.770 63.635 146.795 ;
        RECT 69.995 146.770 70.345 146.795 ;
        RECT 76.705 146.770 77.055 146.795 ;
        RECT 83.415 146.770 83.765 146.795 ;
        RECT 90.125 146.770 90.475 146.795 ;
        RECT 29.240 146.470 30.580 146.770 ;
        RECT 35.950 146.470 37.290 146.770 ;
        RECT 42.660 146.470 44.000 146.770 ;
        RECT 49.370 146.470 50.710 146.770 ;
        RECT 56.080 146.470 57.420 146.770 ;
        RECT 62.790 146.470 64.130 146.770 ;
        RECT 69.500 146.470 70.840 146.770 ;
        RECT 76.210 146.470 77.550 146.770 ;
        RECT 82.920 146.470 84.260 146.770 ;
        RECT 89.630 146.470 90.970 146.770 ;
        RECT 29.735 146.445 30.085 146.470 ;
        RECT 36.445 146.445 36.795 146.470 ;
        RECT 43.155 146.445 43.505 146.470 ;
        RECT 49.865 146.445 50.215 146.470 ;
        RECT 56.575 146.445 56.925 146.470 ;
        RECT 63.285 146.445 63.635 146.470 ;
        RECT 69.995 146.445 70.345 146.470 ;
        RECT 76.705 146.445 77.055 146.470 ;
        RECT 83.415 146.445 83.765 146.470 ;
        RECT 90.125 146.445 90.475 146.470 ;
        RECT 26.730 146.020 27.080 146.045 ;
        RECT 33.440 146.020 33.790 146.045 ;
        RECT 39.000 146.020 41.000 146.075 ;
        RECT 44.000 146.020 46.000 146.075 ;
        RECT 46.860 146.020 47.210 146.045 ;
        RECT 49.000 146.020 51.000 146.075 ;
        RECT 65.000 146.045 67.000 146.075 ;
        RECT 53.570 146.020 53.920 146.045 ;
        RECT 60.280 146.020 60.630 146.045 ;
        RECT 65.000 146.020 67.340 146.045 ;
        RECT 70.000 146.020 72.000 146.075 ;
        RECT 73.700 146.020 74.050 146.045 ;
        RECT 75.000 146.020 77.000 146.075 ;
        RECT 80.410 146.020 80.760 146.045 ;
        RECT 87.120 146.020 87.470 146.045 ;
        RECT 26.730 145.720 93.100 146.020 ;
        RECT 26.730 145.695 27.080 145.720 ;
        RECT 33.440 145.695 33.790 145.720 ;
        RECT 39.000 145.665 41.000 145.720 ;
        RECT 44.000 145.665 46.000 145.720 ;
        RECT 46.860 145.695 47.210 145.720 ;
        RECT 49.000 145.665 51.000 145.720 ;
        RECT 53.570 145.695 53.920 145.720 ;
        RECT 60.280 145.695 60.630 145.720 ;
        RECT 65.000 145.695 67.340 145.720 ;
        RECT 65.000 145.665 67.000 145.695 ;
        RECT 70.000 145.665 72.000 145.720 ;
        RECT 73.700 145.695 74.050 145.720 ;
        RECT 75.000 145.665 77.000 145.720 ;
        RECT 80.410 145.695 80.760 145.720 ;
        RECT 87.120 145.695 87.470 145.720 ;
        RECT 32.390 144.520 32.740 144.545 ;
        RECT 39.000 144.520 41.000 144.575 ;
        RECT 44.000 144.545 46.000 144.575 ;
        RECT 44.000 144.520 46.160 144.545 ;
        RECT 49.000 144.520 51.000 144.575 ;
        RECT 52.520 144.520 52.870 144.545 ;
        RECT 59.230 144.520 59.580 144.545 ;
        RECT 65.000 144.520 67.000 144.575 ;
        RECT 70.000 144.520 72.000 144.575 ;
        RECT 72.650 144.520 73.000 144.545 ;
        RECT 75.000 144.520 77.000 144.575 ;
        RECT 79.360 144.520 79.710 144.545 ;
        RECT 86.070 144.520 86.420 144.545 ;
        RECT 92.780 144.520 93.130 144.545 ;
        RECT 26.760 144.220 93.130 144.520 ;
        RECT 32.390 144.195 32.740 144.220 ;
        RECT 39.000 144.165 41.000 144.220 ;
        RECT 44.000 144.195 46.160 144.220 ;
        RECT 44.000 144.165 46.000 144.195 ;
        RECT 49.000 144.165 51.000 144.220 ;
        RECT 52.520 144.195 52.870 144.220 ;
        RECT 59.230 144.195 59.580 144.220 ;
        RECT 65.000 144.165 67.000 144.220 ;
        RECT 70.000 144.165 72.000 144.220 ;
        RECT 72.650 144.195 73.000 144.220 ;
        RECT 75.000 144.165 77.000 144.220 ;
        RECT 79.360 144.195 79.710 144.220 ;
        RECT 86.070 144.195 86.420 144.220 ;
        RECT 92.780 144.195 93.130 144.220 ;
        RECT 26.730 143.020 27.080 143.045 ;
        RECT 33.440 143.020 33.790 143.045 ;
        RECT 39.000 143.020 41.000 143.075 ;
        RECT 44.000 143.020 46.000 143.075 ;
        RECT 46.860 143.020 47.210 143.045 ;
        RECT 49.000 143.020 51.000 143.075 ;
        RECT 65.000 143.045 67.000 143.075 ;
        RECT 53.570 143.020 53.920 143.045 ;
        RECT 60.280 143.020 60.630 143.045 ;
        RECT 65.000 143.020 67.340 143.045 ;
        RECT 70.000 143.020 72.000 143.075 ;
        RECT 73.700 143.020 74.050 143.045 ;
        RECT 75.000 143.020 77.000 143.075 ;
        RECT 80.410 143.020 80.760 143.045 ;
        RECT 87.120 143.020 87.470 143.045 ;
        RECT 26.730 142.720 93.100 143.020 ;
        RECT 26.730 142.695 27.080 142.720 ;
        RECT 33.440 142.695 33.790 142.720 ;
        RECT 39.000 142.665 41.000 142.720 ;
        RECT 44.000 142.665 46.000 142.720 ;
        RECT 46.860 142.695 47.210 142.720 ;
        RECT 49.000 142.665 51.000 142.720 ;
        RECT 53.570 142.695 53.920 142.720 ;
        RECT 60.280 142.695 60.630 142.720 ;
        RECT 65.000 142.695 67.340 142.720 ;
        RECT 65.000 142.665 67.000 142.695 ;
        RECT 70.000 142.665 72.000 142.720 ;
        RECT 73.700 142.695 74.050 142.720 ;
        RECT 75.000 142.665 77.000 142.720 ;
        RECT 80.410 142.695 80.760 142.720 ;
        RECT 87.120 142.695 87.470 142.720 ;
        RECT 26.250 142.270 26.600 142.295 ;
        RECT 29.735 142.270 30.085 142.295 ;
        RECT 32.960 142.270 33.310 142.295 ;
        RECT 36.445 142.270 36.795 142.295 ;
        RECT 39.670 142.270 40.020 142.295 ;
        RECT 43.155 142.270 43.505 142.295 ;
        RECT 46.380 142.270 46.730 142.295 ;
        RECT 49.865 142.270 50.215 142.295 ;
        RECT 53.090 142.270 53.440 142.295 ;
        RECT 56.575 142.270 56.925 142.295 ;
        RECT 59.800 142.270 60.150 142.295 ;
        RECT 63.285 142.270 63.635 142.295 ;
        RECT 66.510 142.270 66.860 142.295 ;
        RECT 69.995 142.270 70.345 142.295 ;
        RECT 73.220 142.270 73.570 142.295 ;
        RECT 76.705 142.270 77.055 142.295 ;
        RECT 79.930 142.270 80.280 142.295 ;
        RECT 83.415 142.270 83.765 142.295 ;
        RECT 86.640 142.270 86.990 142.295 ;
        RECT 90.125 142.270 90.475 142.295 ;
        RECT 26.250 141.970 30.580 142.270 ;
        RECT 32.960 141.970 37.290 142.270 ;
        RECT 39.670 141.970 44.000 142.270 ;
        RECT 46.380 141.970 50.710 142.270 ;
        RECT 53.090 141.970 57.420 142.270 ;
        RECT 59.800 141.970 64.130 142.270 ;
        RECT 66.510 141.970 70.840 142.270 ;
        RECT 73.220 141.970 77.550 142.270 ;
        RECT 79.930 141.970 84.260 142.270 ;
        RECT 86.640 141.970 90.970 142.270 ;
        RECT 26.250 141.945 26.600 141.970 ;
        RECT 29.735 141.945 30.085 141.970 ;
        RECT 32.960 141.945 33.310 141.970 ;
        RECT 36.445 141.945 36.795 141.970 ;
        RECT 39.670 141.945 40.020 141.970 ;
        RECT 43.155 141.945 43.505 141.970 ;
        RECT 46.380 141.945 46.730 141.970 ;
        RECT 49.865 141.945 50.215 141.970 ;
        RECT 53.090 141.945 53.440 141.970 ;
        RECT 56.575 141.945 56.925 141.970 ;
        RECT 59.800 141.945 60.150 141.970 ;
        RECT 63.285 141.945 63.635 141.970 ;
        RECT 66.510 141.945 66.860 141.970 ;
        RECT 69.995 141.945 70.345 141.970 ;
        RECT 73.220 141.945 73.570 141.970 ;
        RECT 76.705 141.945 77.055 141.970 ;
        RECT 79.930 141.945 80.280 141.970 ;
        RECT 83.415 141.945 83.765 141.970 ;
        RECT 86.640 141.945 86.990 141.970 ;
        RECT 90.125 141.945 90.475 141.970 ;
        RECT 32.390 141.520 32.740 141.545 ;
        RECT 39.000 141.520 41.000 141.575 ;
        RECT 44.000 141.545 46.000 141.575 ;
        RECT 44.000 141.520 46.160 141.545 ;
        RECT 49.000 141.520 51.000 141.575 ;
        RECT 52.520 141.520 52.870 141.545 ;
        RECT 59.230 141.520 59.580 141.545 ;
        RECT 65.000 141.520 67.000 141.575 ;
        RECT 70.000 141.520 72.000 141.575 ;
        RECT 72.650 141.520 73.000 141.545 ;
        RECT 75.000 141.520 77.000 141.575 ;
        RECT 79.360 141.520 79.710 141.545 ;
        RECT 86.070 141.520 86.420 141.545 ;
        RECT 92.780 141.520 93.130 141.545 ;
        RECT 26.760 141.220 93.130 141.520 ;
        RECT 32.390 141.195 32.740 141.220 ;
        RECT 39.000 141.165 41.000 141.220 ;
        RECT 44.000 141.195 46.160 141.220 ;
        RECT 44.000 141.165 46.000 141.195 ;
        RECT 49.000 141.165 51.000 141.220 ;
        RECT 52.520 141.195 52.870 141.220 ;
        RECT 59.230 141.195 59.580 141.220 ;
        RECT 65.000 141.165 67.000 141.220 ;
        RECT 70.000 141.165 72.000 141.220 ;
        RECT 72.650 141.195 73.000 141.220 ;
        RECT 75.000 141.165 77.000 141.220 ;
        RECT 79.360 141.195 79.710 141.220 ;
        RECT 86.070 141.195 86.420 141.220 ;
        RECT 92.780 141.195 93.130 141.220 ;
        RECT 26.730 140.020 27.080 140.045 ;
        RECT 33.440 140.020 33.790 140.045 ;
        RECT 39.000 140.020 41.000 140.075 ;
        RECT 44.000 140.020 46.000 140.075 ;
        RECT 46.860 140.020 47.210 140.045 ;
        RECT 49.000 140.020 51.000 140.075 ;
        RECT 65.000 140.045 67.000 140.075 ;
        RECT 53.570 140.020 53.920 140.045 ;
        RECT 60.280 140.020 60.630 140.045 ;
        RECT 65.000 140.020 67.340 140.045 ;
        RECT 70.000 140.020 72.000 140.075 ;
        RECT 73.700 140.020 74.050 140.045 ;
        RECT 75.000 140.020 77.000 140.075 ;
        RECT 80.410 140.020 80.760 140.045 ;
        RECT 87.120 140.020 87.470 140.045 ;
        RECT 26.730 139.720 93.100 140.020 ;
        RECT 26.730 139.695 27.080 139.720 ;
        RECT 33.440 139.695 33.790 139.720 ;
        RECT 39.000 139.665 41.000 139.720 ;
        RECT 44.000 139.665 46.000 139.720 ;
        RECT 46.860 139.695 47.210 139.720 ;
        RECT 49.000 139.665 51.000 139.720 ;
        RECT 53.570 139.695 53.920 139.720 ;
        RECT 60.280 139.695 60.630 139.720 ;
        RECT 65.000 139.695 67.340 139.720 ;
        RECT 65.000 139.665 67.000 139.695 ;
        RECT 70.000 139.665 72.000 139.720 ;
        RECT 73.700 139.695 74.050 139.720 ;
        RECT 75.000 139.665 77.000 139.720 ;
        RECT 80.410 139.695 80.760 139.720 ;
        RECT 87.120 139.695 87.470 139.720 ;
        RECT 31.540 139.270 31.890 139.295 ;
        RECT 35.550 139.270 35.900 139.295 ;
        RECT 31.540 138.970 35.900 139.270 ;
        RECT 31.540 138.945 31.890 138.970 ;
        RECT 35.550 138.945 35.900 138.970 ;
        RECT 44.960 139.270 45.310 139.295 ;
        RECT 48.970 139.270 49.320 139.295 ;
        RECT 44.960 138.970 49.320 139.270 ;
        RECT 44.960 138.945 45.310 138.970 ;
        RECT 48.970 138.945 49.320 138.970 ;
        RECT 58.380 139.270 58.730 139.295 ;
        RECT 62.390 139.270 62.740 139.295 ;
        RECT 58.380 138.970 62.740 139.270 ;
        RECT 58.380 138.945 58.730 138.970 ;
        RECT 62.390 138.945 62.740 138.970 ;
        RECT 71.800 139.270 72.150 139.295 ;
        RECT 75.810 139.270 76.160 139.295 ;
        RECT 71.800 138.970 76.160 139.270 ;
        RECT 71.800 138.945 72.150 138.970 ;
        RECT 75.810 138.945 76.160 138.970 ;
        RECT 85.220 139.270 85.570 139.295 ;
        RECT 89.230 139.270 89.580 139.295 ;
        RECT 85.220 138.970 89.580 139.270 ;
        RECT 85.220 138.945 85.570 138.970 ;
        RECT 89.230 138.945 89.580 138.970 ;
        RECT 32.390 138.520 32.740 138.545 ;
        RECT 39.000 138.520 41.000 138.575 ;
        RECT 44.000 138.545 46.000 138.575 ;
        RECT 44.000 138.520 46.160 138.545 ;
        RECT 49.000 138.520 51.000 138.575 ;
        RECT 52.520 138.520 52.870 138.545 ;
        RECT 59.230 138.520 59.580 138.545 ;
        RECT 65.000 138.520 67.000 138.575 ;
        RECT 70.000 138.520 72.000 138.575 ;
        RECT 72.650 138.520 73.000 138.545 ;
        RECT 75.000 138.520 77.000 138.575 ;
        RECT 79.360 138.520 79.710 138.545 ;
        RECT 86.070 138.520 86.420 138.545 ;
        RECT 92.780 138.520 93.130 138.545 ;
        RECT 26.760 138.220 93.130 138.520 ;
        RECT 32.390 138.195 32.740 138.220 ;
        RECT 39.000 138.165 41.000 138.220 ;
        RECT 44.000 138.195 46.160 138.220 ;
        RECT 44.000 138.165 46.000 138.195 ;
        RECT 49.000 138.165 51.000 138.220 ;
        RECT 52.520 138.195 52.870 138.220 ;
        RECT 59.230 138.195 59.580 138.220 ;
        RECT 65.000 138.165 67.000 138.220 ;
        RECT 70.000 138.165 72.000 138.220 ;
        RECT 72.650 138.195 73.000 138.220 ;
        RECT 75.000 138.165 77.000 138.220 ;
        RECT 79.360 138.195 79.710 138.220 ;
        RECT 86.070 138.195 86.420 138.220 ;
        RECT 92.780 138.195 93.130 138.220 ;
        RECT 28.000 137.770 28.350 137.795 ;
        RECT 34.710 137.770 35.060 137.795 ;
        RECT 28.000 137.470 35.060 137.770 ;
        RECT 28.000 137.445 28.350 137.470 ;
        RECT 34.710 137.445 35.060 137.470 ;
        RECT 41.420 137.770 41.770 137.795 ;
        RECT 48.130 137.770 48.480 137.795 ;
        RECT 41.420 137.470 48.480 137.770 ;
        RECT 41.420 137.445 41.770 137.470 ;
        RECT 48.130 137.445 48.480 137.470 ;
        RECT 54.840 137.770 55.190 137.795 ;
        RECT 61.550 137.770 61.900 137.795 ;
        RECT 54.840 137.470 61.900 137.770 ;
        RECT 54.840 137.445 55.190 137.470 ;
        RECT 61.550 137.445 61.900 137.470 ;
        RECT 68.260 137.770 68.610 137.795 ;
        RECT 74.970 137.770 75.320 137.795 ;
        RECT 68.260 137.470 75.320 137.770 ;
        RECT 68.260 137.445 68.610 137.470 ;
        RECT 74.970 137.445 75.320 137.470 ;
        RECT 81.680 137.770 82.030 137.795 ;
        RECT 88.390 137.770 88.740 137.795 ;
        RECT 81.680 137.470 88.740 137.770 ;
        RECT 81.680 137.445 82.030 137.470 ;
        RECT 88.390 137.445 88.740 137.470 ;
        RECT 26.730 137.020 27.080 137.045 ;
        RECT 33.440 137.020 33.790 137.045 ;
        RECT 39.000 137.020 41.000 137.075 ;
        RECT 44.000 137.020 46.000 137.075 ;
        RECT 46.860 137.020 47.210 137.045 ;
        RECT 49.000 137.020 51.000 137.075 ;
        RECT 65.000 137.045 67.000 137.075 ;
        RECT 53.570 137.020 53.920 137.045 ;
        RECT 60.280 137.020 60.630 137.045 ;
        RECT 65.000 137.020 67.340 137.045 ;
        RECT 70.000 137.020 72.000 137.075 ;
        RECT 73.700 137.020 74.050 137.045 ;
        RECT 75.000 137.020 77.000 137.075 ;
        RECT 80.410 137.020 80.760 137.045 ;
        RECT 87.120 137.020 87.470 137.045 ;
        RECT 26.730 136.720 93.100 137.020 ;
        RECT 26.730 136.695 27.080 136.720 ;
        RECT 33.440 136.695 33.790 136.720 ;
        RECT 39.000 136.665 41.000 136.720 ;
        RECT 44.000 136.665 46.000 136.720 ;
        RECT 46.860 136.695 47.210 136.720 ;
        RECT 49.000 136.665 51.000 136.720 ;
        RECT 53.570 136.695 53.920 136.720 ;
        RECT 60.280 136.695 60.630 136.720 ;
        RECT 65.000 136.695 67.340 136.720 ;
        RECT 65.000 136.665 67.000 136.695 ;
        RECT 70.000 136.665 72.000 136.720 ;
        RECT 73.700 136.695 74.050 136.720 ;
        RECT 75.000 136.665 77.000 136.720 ;
        RECT 80.410 136.695 80.760 136.720 ;
        RECT 87.120 136.695 87.470 136.720 ;
        RECT 28.420 136.270 28.770 136.295 ;
        RECT 35.130 136.270 35.480 136.295 ;
        RECT 28.420 135.970 35.480 136.270 ;
        RECT 28.420 135.945 28.770 135.970 ;
        RECT 35.130 135.945 35.480 135.970 ;
        RECT 41.840 136.270 42.190 136.295 ;
        RECT 48.550 136.270 48.900 136.295 ;
        RECT 41.840 135.970 48.900 136.270 ;
        RECT 41.840 135.945 42.190 135.970 ;
        RECT 48.550 135.945 48.900 135.970 ;
        RECT 55.260 136.270 55.610 136.295 ;
        RECT 61.970 136.270 62.320 136.295 ;
        RECT 55.260 135.970 62.320 136.270 ;
        RECT 55.260 135.945 55.610 135.970 ;
        RECT 61.970 135.945 62.320 135.970 ;
        RECT 68.680 136.270 69.030 136.295 ;
        RECT 75.390 136.270 75.740 136.295 ;
        RECT 68.680 135.970 75.740 136.270 ;
        RECT 68.680 135.945 69.030 135.970 ;
        RECT 75.390 135.945 75.740 135.970 ;
        RECT 82.100 136.270 82.450 136.295 ;
        RECT 88.810 136.270 89.160 136.295 ;
        RECT 82.100 135.970 89.160 136.270 ;
        RECT 82.100 135.945 82.450 135.970 ;
        RECT 88.810 135.945 89.160 135.970 ;
        RECT 32.390 135.520 32.740 135.545 ;
        RECT 39.000 135.520 41.000 135.575 ;
        RECT 44.000 135.545 46.000 135.575 ;
        RECT 44.000 135.520 46.160 135.545 ;
        RECT 49.000 135.520 51.000 135.575 ;
        RECT 52.520 135.520 52.870 135.545 ;
        RECT 59.230 135.520 59.580 135.545 ;
        RECT 65.000 135.520 67.000 135.575 ;
        RECT 70.000 135.520 72.000 135.575 ;
        RECT 72.650 135.520 73.000 135.545 ;
        RECT 75.000 135.520 77.000 135.575 ;
        RECT 79.360 135.520 79.710 135.545 ;
        RECT 86.070 135.520 86.420 135.545 ;
        RECT 92.780 135.520 93.130 135.545 ;
        RECT 26.760 135.220 93.130 135.520 ;
        RECT 32.390 135.195 32.740 135.220 ;
        RECT 39.000 135.165 41.000 135.220 ;
        RECT 44.000 135.195 46.160 135.220 ;
        RECT 44.000 135.165 46.000 135.195 ;
        RECT 49.000 135.165 51.000 135.220 ;
        RECT 52.520 135.195 52.870 135.220 ;
        RECT 59.230 135.195 59.580 135.220 ;
        RECT 65.000 135.165 67.000 135.220 ;
        RECT 70.000 135.165 72.000 135.220 ;
        RECT 72.650 135.195 73.000 135.220 ;
        RECT 75.000 135.165 77.000 135.220 ;
        RECT 79.360 135.195 79.710 135.220 ;
        RECT 86.070 135.195 86.420 135.220 ;
        RECT 92.780 135.195 93.130 135.220 ;
        RECT 27.580 134.770 27.930 134.795 ;
        RECT 34.290 134.770 34.640 134.795 ;
        RECT 27.580 134.470 34.640 134.770 ;
        RECT 27.580 134.445 27.930 134.470 ;
        RECT 34.290 134.445 34.640 134.470 ;
        RECT 41.000 134.770 41.350 134.795 ;
        RECT 47.710 134.770 48.060 134.795 ;
        RECT 41.000 134.470 48.060 134.770 ;
        RECT 41.000 134.445 41.350 134.470 ;
        RECT 47.710 134.445 48.060 134.470 ;
        RECT 54.420 134.770 54.770 134.795 ;
        RECT 61.130 134.770 61.480 134.795 ;
        RECT 54.420 134.470 61.480 134.770 ;
        RECT 54.420 134.445 54.770 134.470 ;
        RECT 61.130 134.445 61.480 134.470 ;
        RECT 67.840 134.770 68.190 134.795 ;
        RECT 74.550 134.770 74.900 134.795 ;
        RECT 67.840 134.470 74.900 134.770 ;
        RECT 67.840 134.445 68.190 134.470 ;
        RECT 74.550 134.445 74.900 134.470 ;
        RECT 81.260 134.770 81.610 134.795 ;
        RECT 87.970 134.770 88.320 134.795 ;
        RECT 81.260 134.470 88.320 134.770 ;
        RECT 81.260 134.445 81.610 134.470 ;
        RECT 87.970 134.445 88.320 134.470 ;
        RECT 26.730 134.020 27.080 134.045 ;
        RECT 33.440 134.020 33.790 134.045 ;
        RECT 39.000 134.020 41.000 134.075 ;
        RECT 44.000 134.020 46.000 134.075 ;
        RECT 46.860 134.020 47.210 134.045 ;
        RECT 49.000 134.020 51.000 134.075 ;
        RECT 65.000 134.045 67.000 134.075 ;
        RECT 53.570 134.020 53.920 134.045 ;
        RECT 60.280 134.020 60.630 134.045 ;
        RECT 65.000 134.020 67.340 134.045 ;
        RECT 70.000 134.020 72.000 134.075 ;
        RECT 73.700 134.020 74.050 134.045 ;
        RECT 75.000 134.020 77.000 134.075 ;
        RECT 80.410 134.020 80.760 134.045 ;
        RECT 87.120 134.020 87.470 134.045 ;
        RECT 26.730 133.720 93.100 134.020 ;
        RECT 26.730 133.695 27.080 133.720 ;
        RECT 33.440 133.695 33.790 133.720 ;
        RECT 39.000 133.665 41.000 133.720 ;
        RECT 44.000 133.665 46.000 133.720 ;
        RECT 46.860 133.695 47.210 133.720 ;
        RECT 49.000 133.665 51.000 133.720 ;
        RECT 53.570 133.695 53.920 133.720 ;
        RECT 60.280 133.695 60.630 133.720 ;
        RECT 65.000 133.695 67.340 133.720 ;
        RECT 65.000 133.665 67.000 133.695 ;
        RECT 70.000 133.665 72.000 133.720 ;
        RECT 73.700 133.695 74.050 133.720 ;
        RECT 75.000 133.665 77.000 133.720 ;
        RECT 80.410 133.695 80.760 133.720 ;
        RECT 87.120 133.695 87.470 133.720 ;
        RECT 107.000 123.000 109.000 123.030 ;
        RECT 16.000 121.000 119.000 123.000 ;
        RECT 107.000 120.970 109.000 121.000 ;
        RECT 16.000 118.000 18.000 118.030 ;
        RECT 44.000 118.000 46.000 118.030 ;
        RECT 16.000 116.000 119.000 118.000 ;
        RECT 16.000 115.970 18.000 116.000 ;
        RECT 44.000 115.970 46.000 116.000 ;
        RECT 49.000 113.000 51.000 113.030 ;
        RECT 75.000 113.000 77.000 113.030 ;
        RECT 117.000 113.000 119.000 113.030 ;
        RECT 16.000 111.000 119.000 113.000 ;
        RECT 49.000 110.970 51.000 111.000 ;
        RECT 75.000 110.970 77.000 111.000 ;
        RECT 117.000 110.970 119.000 111.000 ;
        RECT 39.000 103.010 41.000 103.040 ;
        RECT 33.775 102.010 46.075 103.010 ;
        RECT 33.775 100.840 34.075 102.010 ;
        RECT 36.775 100.840 37.075 102.010 ;
        RECT 39.000 101.980 41.000 102.010 ;
        RECT 39.775 100.840 40.075 101.980 ;
        RECT 42.000 100.970 42.350 101.320 ;
        RECT 33.750 100.490 34.100 100.840 ;
        RECT 33.775 94.130 34.075 100.490 ;
        RECT 34.500 99.640 34.850 99.990 ;
        RECT 33.750 93.780 34.100 94.130 ;
        RECT 33.775 87.420 34.075 93.780 ;
        RECT 34.525 93.280 34.825 99.640 ;
        RECT 35.275 95.180 35.575 100.810 ;
        RECT 36.750 100.490 37.100 100.840 ;
        RECT 39.750 100.810 40.100 100.840 ;
        RECT 36.000 98.800 36.350 99.150 ;
        RECT 35.250 94.830 35.600 95.180 ;
        RECT 34.500 92.930 34.850 93.280 ;
        RECT 35.275 88.470 35.575 94.830 ;
        RECT 36.025 92.440 36.325 98.800 ;
        RECT 36.775 94.130 37.075 100.490 ;
        RECT 37.500 99.220 37.850 99.570 ;
        RECT 36.750 93.780 37.100 94.130 ;
        RECT 36.000 92.090 36.350 92.440 ;
        RECT 35.250 88.120 35.600 88.470 ;
        RECT 33.750 87.070 34.100 87.420 ;
        RECT 33.775 80.710 34.075 87.070 ;
        RECT 34.500 86.220 34.850 86.570 ;
        RECT 33.750 80.360 34.100 80.710 ;
        RECT 33.775 74.000 34.075 80.360 ;
        RECT 34.525 79.860 34.825 86.220 ;
        RECT 35.275 81.760 35.575 88.120 ;
        RECT 36.775 87.420 37.075 93.780 ;
        RECT 37.525 92.860 37.825 99.220 ;
        RECT 38.275 95.180 38.575 100.810 ;
        RECT 39.000 95.680 39.350 96.030 ;
        RECT 38.250 94.830 38.600 95.180 ;
        RECT 37.500 92.510 37.850 92.860 ;
        RECT 38.275 88.470 38.575 94.830 ;
        RECT 39.025 92.020 39.325 95.680 ;
        RECT 39.000 91.670 39.350 92.020 ;
        RECT 38.250 88.120 38.600 88.470 ;
        RECT 36.750 87.070 37.100 87.420 ;
        RECT 36.000 85.380 36.350 85.730 ;
        RECT 35.250 81.410 35.600 81.760 ;
        RECT 34.500 79.510 34.850 79.860 ;
        RECT 35.275 75.050 35.575 81.410 ;
        RECT 36.025 79.020 36.325 85.380 ;
        RECT 36.775 80.710 37.075 87.070 ;
        RECT 37.500 85.800 37.850 86.150 ;
        RECT 36.750 80.360 37.100 80.710 ;
        RECT 36.000 78.670 36.350 79.020 ;
        RECT 35.250 74.700 35.600 75.050 ;
        RECT 33.750 73.650 34.100 74.000 ;
        RECT 33.775 67.290 34.075 73.650 ;
        RECT 34.500 72.800 34.850 73.150 ;
        RECT 33.750 66.940 34.100 67.290 ;
        RECT 33.775 60.580 34.075 66.940 ;
        RECT 34.525 66.440 34.825 72.800 ;
        RECT 35.275 68.340 35.575 74.700 ;
        RECT 36.775 74.000 37.075 80.360 ;
        RECT 37.525 79.440 37.825 85.800 ;
        RECT 38.275 81.760 38.575 88.120 ;
        RECT 39.000 82.260 39.350 82.610 ;
        RECT 38.250 81.410 38.600 81.760 ;
        RECT 37.500 79.090 37.850 79.440 ;
        RECT 38.275 75.050 38.575 81.410 ;
        RECT 39.025 78.600 39.325 82.260 ;
        RECT 39.000 78.250 39.350 78.600 ;
        RECT 38.250 74.700 38.600 75.050 ;
        RECT 36.750 73.650 37.100 74.000 ;
        RECT 36.000 71.960 36.350 72.310 ;
        RECT 35.250 67.990 35.600 68.340 ;
        RECT 34.500 66.090 34.850 66.440 ;
        RECT 35.275 61.630 35.575 67.990 ;
        RECT 36.025 65.600 36.325 71.960 ;
        RECT 36.775 67.290 37.075 73.650 ;
        RECT 37.500 72.380 37.850 72.730 ;
        RECT 36.750 66.940 37.100 67.290 ;
        RECT 36.000 65.250 36.350 65.600 ;
        RECT 35.250 61.280 35.600 61.630 ;
        RECT 33.750 60.230 34.100 60.580 ;
        RECT 33.775 53.870 34.075 60.230 ;
        RECT 34.500 59.380 34.850 59.730 ;
        RECT 33.750 53.520 34.100 53.870 ;
        RECT 33.775 47.160 34.075 53.520 ;
        RECT 34.525 53.020 34.825 59.380 ;
        RECT 35.275 54.920 35.575 61.280 ;
        RECT 36.775 60.580 37.075 66.940 ;
        RECT 37.525 66.020 37.825 72.380 ;
        RECT 38.275 68.340 38.575 74.700 ;
        RECT 39.000 68.840 39.350 69.190 ;
        RECT 38.250 67.990 38.600 68.340 ;
        RECT 37.500 65.670 37.850 66.020 ;
        RECT 38.275 61.630 38.575 67.990 ;
        RECT 39.025 65.180 39.325 68.840 ;
        RECT 39.000 64.830 39.350 65.180 ;
        RECT 38.250 61.280 38.600 61.630 ;
        RECT 36.750 60.230 37.100 60.580 ;
        RECT 36.000 58.540 36.350 58.890 ;
        RECT 35.250 54.570 35.600 54.920 ;
        RECT 34.500 52.670 34.850 53.020 ;
        RECT 35.275 48.210 35.575 54.570 ;
        RECT 36.025 52.180 36.325 58.540 ;
        RECT 36.775 53.870 37.075 60.230 ;
        RECT 37.500 58.960 37.850 59.310 ;
        RECT 36.750 53.520 37.100 53.870 ;
        RECT 36.000 51.830 36.350 52.180 ;
        RECT 35.250 47.860 35.600 48.210 ;
        RECT 33.750 46.810 34.100 47.160 ;
        RECT 33.775 40.450 34.075 46.810 ;
        RECT 34.500 45.960 34.850 46.310 ;
        RECT 33.750 40.100 34.100 40.450 ;
        RECT 33.775 34.470 34.075 40.100 ;
        RECT 34.525 39.600 34.825 45.960 ;
        RECT 35.275 41.500 35.575 47.860 ;
        RECT 36.775 47.160 37.075 53.520 ;
        RECT 37.525 52.600 37.825 58.960 ;
        RECT 38.275 54.920 38.575 61.280 ;
        RECT 39.000 55.420 39.350 55.770 ;
        RECT 38.250 54.570 38.600 54.920 ;
        RECT 37.500 52.250 37.850 52.600 ;
        RECT 38.275 48.210 38.575 54.570 ;
        RECT 39.025 51.760 39.325 55.420 ;
        RECT 39.000 51.410 39.350 51.760 ;
        RECT 38.250 47.860 38.600 48.210 ;
        RECT 36.750 46.810 37.100 47.160 ;
        RECT 36.000 45.120 36.350 45.470 ;
        RECT 35.250 41.150 35.600 41.500 ;
        RECT 34.500 39.250 34.850 39.600 ;
        RECT 35.275 34.790 35.575 41.150 ;
        RECT 36.025 38.760 36.325 45.120 ;
        RECT 36.775 40.450 37.075 46.810 ;
        RECT 37.500 45.540 37.850 45.890 ;
        RECT 36.750 40.100 37.100 40.450 ;
        RECT 36.000 38.410 36.350 38.760 ;
        RECT 35.250 34.440 35.600 34.790 ;
        RECT 36.775 34.470 37.075 40.100 ;
        RECT 37.525 39.180 37.825 45.540 ;
        RECT 38.275 41.500 38.575 47.860 ;
        RECT 39.000 42.000 39.350 42.350 ;
        RECT 38.250 41.150 38.600 41.500 ;
        RECT 37.500 38.830 37.850 39.180 ;
        RECT 38.275 34.790 38.575 41.150 ;
        RECT 39.025 38.340 39.325 42.000 ;
        RECT 39.000 37.990 39.350 38.340 ;
        RECT 38.250 34.440 38.600 34.790 ;
        RECT 39.735 34.470 40.115 100.810 ;
        RECT 41.275 95.180 41.575 100.810 ;
        RECT 42.025 97.835 42.325 100.970 ;
        RECT 42.775 100.840 43.075 102.010 ;
        RECT 45.775 100.840 46.075 102.010 ;
        RECT 42.750 100.490 43.100 100.840 ;
        RECT 42.000 97.485 42.350 97.835 ;
        RECT 42.025 96.990 42.325 97.485 ;
        RECT 41.250 94.830 41.600 95.180 ;
        RECT 41.275 88.470 41.575 94.830 ;
        RECT 42.000 94.260 42.350 94.610 ;
        RECT 42.025 91.125 42.325 94.260 ;
        RECT 42.775 94.130 43.075 100.490 ;
        RECT 42.750 93.780 43.100 94.130 ;
        RECT 42.000 90.775 42.350 91.125 ;
        RECT 42.025 90.280 42.325 90.775 ;
        RECT 41.250 88.120 41.600 88.470 ;
        RECT 41.275 81.760 41.575 88.120 ;
        RECT 42.000 87.550 42.350 87.900 ;
        RECT 42.025 84.415 42.325 87.550 ;
        RECT 42.775 87.420 43.075 93.780 ;
        RECT 42.750 87.070 43.100 87.420 ;
        RECT 42.000 84.065 42.350 84.415 ;
        RECT 42.025 83.570 42.325 84.065 ;
        RECT 41.250 81.410 41.600 81.760 ;
        RECT 41.275 75.050 41.575 81.410 ;
        RECT 42.000 80.840 42.350 81.190 ;
        RECT 42.025 77.705 42.325 80.840 ;
        RECT 42.775 80.710 43.075 87.070 ;
        RECT 42.750 80.360 43.100 80.710 ;
        RECT 42.000 77.355 42.350 77.705 ;
        RECT 42.025 76.860 42.325 77.355 ;
        RECT 41.250 74.700 41.600 75.050 ;
        RECT 41.275 68.340 41.575 74.700 ;
        RECT 42.000 74.130 42.350 74.480 ;
        RECT 42.025 70.995 42.325 74.130 ;
        RECT 42.775 74.000 43.075 80.360 ;
        RECT 42.750 73.650 43.100 74.000 ;
        RECT 42.000 70.645 42.350 70.995 ;
        RECT 42.025 70.150 42.325 70.645 ;
        RECT 41.250 67.990 41.600 68.340 ;
        RECT 41.275 61.630 41.575 67.990 ;
        RECT 42.000 67.420 42.350 67.770 ;
        RECT 42.025 64.285 42.325 67.420 ;
        RECT 42.775 67.290 43.075 73.650 ;
        RECT 42.750 66.940 43.100 67.290 ;
        RECT 42.000 63.935 42.350 64.285 ;
        RECT 42.025 63.440 42.325 63.935 ;
        RECT 41.250 61.280 41.600 61.630 ;
        RECT 41.275 54.920 41.575 61.280 ;
        RECT 42.000 60.710 42.350 61.060 ;
        RECT 42.025 57.575 42.325 60.710 ;
        RECT 42.775 60.580 43.075 66.940 ;
        RECT 42.750 60.230 43.100 60.580 ;
        RECT 42.000 57.225 42.350 57.575 ;
        RECT 42.025 56.730 42.325 57.225 ;
        RECT 41.250 54.570 41.600 54.920 ;
        RECT 41.275 48.210 41.575 54.570 ;
        RECT 42.000 54.000 42.350 54.350 ;
        RECT 42.025 50.865 42.325 54.000 ;
        RECT 42.775 53.870 43.075 60.230 ;
        RECT 42.750 53.520 43.100 53.870 ;
        RECT 42.000 50.515 42.350 50.865 ;
        RECT 42.025 50.020 42.325 50.515 ;
        RECT 41.250 47.860 41.600 48.210 ;
        RECT 41.275 41.500 41.575 47.860 ;
        RECT 42.000 47.290 42.350 47.640 ;
        RECT 42.025 44.155 42.325 47.290 ;
        RECT 42.775 47.160 43.075 53.520 ;
        RECT 42.750 46.810 43.100 47.160 ;
        RECT 42.000 43.805 42.350 44.155 ;
        RECT 42.025 43.310 42.325 43.805 ;
        RECT 41.250 41.150 41.600 41.500 ;
        RECT 41.275 34.790 41.575 41.150 ;
        RECT 42.000 40.580 42.350 40.930 ;
        RECT 42.025 37.445 42.325 40.580 ;
        RECT 42.775 40.450 43.075 46.810 ;
        RECT 42.750 40.100 43.100 40.450 ;
        RECT 42.000 37.095 42.350 37.445 ;
        RECT 42.025 36.600 42.325 37.095 ;
        RECT 41.250 34.440 41.600 34.790 ;
        RECT 42.775 34.470 43.075 40.100 ;
        RECT 44.235 34.470 44.615 100.810 ;
        RECT 45.750 100.490 46.100 100.840 ;
        RECT 45.775 94.130 46.075 100.490 ;
        RECT 65.485 98.980 66.515 100.070 ;
        RECT 46.525 97.835 46.825 98.330 ;
        RECT 47.155 98.075 67.070 98.375 ;
        RECT 46.500 97.485 46.850 97.835 ;
        RECT 46.525 96.990 46.825 97.485 ;
        RECT 47.155 94.610 47.455 98.075 ;
        RECT 47.785 97.445 65.690 97.745 ;
        RECT 47.130 94.260 47.480 94.610 ;
        RECT 45.750 93.780 46.100 94.130 ;
        RECT 45.775 87.420 46.075 93.780 ;
        RECT 46.525 91.125 46.825 91.620 ;
        RECT 47.785 91.125 48.085 97.445 ;
        RECT 48.390 97.115 48.740 97.140 ;
        RECT 48.390 96.815 64.310 97.115 ;
        RECT 48.390 96.790 48.740 96.815 ;
        RECT 49.020 96.485 49.370 96.510 ;
        RECT 49.020 96.185 62.930 96.485 ;
        RECT 49.020 96.160 49.370 96.185 ;
        RECT 48.415 95.555 61.550 95.855 ;
        RECT 46.500 90.775 46.850 91.125 ;
        RECT 47.760 90.775 48.110 91.125 ;
        RECT 46.525 90.280 46.825 90.775 ;
        RECT 47.130 90.145 47.480 90.495 ;
        RECT 47.155 87.900 47.455 90.145 ;
        RECT 47.760 89.515 48.110 89.865 ;
        RECT 47.130 87.550 47.480 87.900 ;
        RECT 45.750 87.070 46.100 87.420 ;
        RECT 45.775 80.710 46.075 87.070 ;
        RECT 46.525 84.415 46.825 84.910 ;
        RECT 47.785 84.415 48.085 89.515 ;
        RECT 46.500 84.065 46.850 84.415 ;
        RECT 47.760 84.065 48.110 84.415 ;
        RECT 46.525 83.570 46.825 84.065 ;
        RECT 48.415 81.190 48.715 95.555 ;
        RECT 49.045 94.925 60.170 95.225 ;
        RECT 48.390 80.840 48.740 81.190 ;
        RECT 45.750 80.360 46.100 80.710 ;
        RECT 45.775 74.000 46.075 80.360 ;
        RECT 46.525 77.705 46.825 78.200 ;
        RECT 49.045 77.705 49.345 94.925 ;
        RECT 49.675 94.295 58.790 94.595 ;
        RECT 49.675 90.495 49.975 94.295 ;
        RECT 58.490 93.995 58.790 94.295 ;
        RECT 59.870 93.995 60.170 94.925 ;
        RECT 61.250 93.995 61.550 95.555 ;
        RECT 62.630 93.995 62.930 96.185 ;
        RECT 64.010 93.995 64.310 96.815 ;
        RECT 65.390 93.995 65.690 97.445 ;
        RECT 66.770 93.995 67.070 98.075 ;
        RECT 56.965 93.850 57.555 93.995 ;
        RECT 50.305 93.550 57.555 93.850 ;
        RECT 49.650 90.145 50.000 90.495 ;
        RECT 50.305 89.865 50.605 93.550 ;
        RECT 56.965 93.405 57.555 93.550 ;
        RECT 58.345 93.405 58.935 93.995 ;
        RECT 59.725 93.405 60.315 93.995 ;
        RECT 61.105 93.405 61.695 93.995 ;
        RECT 62.485 93.405 63.075 93.995 ;
        RECT 63.865 93.405 64.455 93.995 ;
        RECT 65.245 93.405 65.835 93.995 ;
        RECT 66.625 93.405 67.215 93.995 ;
        RECT 56.915 92.005 69.850 92.695 ;
        RECT 56.915 92.000 57.215 92.005 ;
        RECT 58.295 92.000 58.595 92.005 ;
        RECT 59.675 92.000 59.975 92.005 ;
        RECT 61.055 92.000 61.355 92.005 ;
        RECT 62.435 92.000 62.735 92.005 ;
        RECT 63.815 92.000 64.115 92.005 ;
        RECT 65.195 92.000 65.495 92.005 ;
        RECT 66.575 92.000 66.875 92.005 ;
        RECT 50.280 89.515 50.630 89.865 ;
        RECT 57.425 89.075 58.115 89.465 ;
        RECT 50.600 88.775 58.115 89.075 ;
        RECT 58.805 88.775 59.495 89.465 ;
        RECT 60.185 88.775 60.875 89.465 ;
        RECT 61.565 88.775 62.255 89.465 ;
        RECT 62.945 88.775 63.635 89.465 ;
        RECT 64.325 88.775 65.015 89.465 ;
        RECT 65.705 88.775 66.395 89.465 ;
        RECT 67.085 88.775 67.775 89.465 ;
        RECT 50.600 85.765 50.900 88.775 ;
        RECT 58.805 88.450 59.105 88.775 ;
        RECT 52.260 88.150 59.105 88.450 ;
        RECT 52.260 85.765 52.560 88.150 ;
        RECT 60.185 87.825 60.485 88.775 ;
        RECT 53.920 87.525 60.485 87.825 ;
        RECT 53.920 85.765 54.220 87.525 ;
        RECT 61.565 87.200 61.865 88.775 ;
        RECT 55.580 86.900 61.865 87.200 ;
        RECT 55.580 85.765 55.880 86.900 ;
        RECT 62.945 86.575 63.245 88.775 ;
        RECT 57.240 86.275 63.245 86.575 ;
        RECT 57.240 85.765 57.540 86.275 ;
        RECT 64.325 85.950 64.625 88.775 ;
        RECT 58.900 85.765 64.625 85.950 ;
        RECT 50.575 85.415 50.925 85.765 ;
        RECT 52.235 85.415 52.585 85.765 ;
        RECT 53.895 85.415 54.245 85.765 ;
        RECT 55.555 85.415 55.905 85.765 ;
        RECT 57.215 85.415 57.565 85.765 ;
        RECT 58.875 85.650 64.625 85.765 ;
        RECT 58.875 85.415 59.225 85.650 ;
        RECT 60.535 85.325 60.885 85.350 ;
        RECT 65.705 85.325 66.005 88.775 ;
        RECT 60.535 85.025 66.005 85.325 ;
        RECT 60.535 85.000 60.885 85.025 ;
        RECT 62.195 84.700 62.545 84.725 ;
        RECT 67.085 84.700 67.385 88.775 ;
        RECT 62.195 84.400 67.385 84.700 ;
        RECT 62.195 84.375 62.545 84.400 ;
        RECT 46.500 77.355 46.850 77.705 ;
        RECT 49.020 77.355 49.370 77.705 ;
        RECT 46.525 76.860 46.825 77.355 ;
        RECT 51.540 74.130 51.890 74.480 ;
        RECT 45.750 73.650 46.100 74.000 ;
        RECT 45.775 67.290 46.075 73.650 ;
        RECT 46.525 70.995 46.825 71.490 ;
        RECT 46.500 70.645 46.850 70.995 ;
        RECT 50.910 70.645 51.260 70.995 ;
        RECT 46.525 70.150 46.825 70.645 ;
        RECT 47.130 67.420 47.480 67.770 ;
        RECT 45.750 66.940 46.100 67.290 ;
        RECT 45.775 60.580 46.075 66.940 ;
        RECT 46.525 64.285 46.825 64.780 ;
        RECT 46.500 63.935 46.850 64.285 ;
        RECT 46.525 63.440 46.825 63.935 ;
        RECT 45.750 60.230 46.100 60.580 ;
        RECT 45.775 53.870 46.075 60.230 ;
        RECT 46.525 57.575 46.825 58.070 ;
        RECT 46.500 57.225 46.850 57.575 ;
        RECT 46.525 56.730 46.825 57.225 ;
        RECT 45.750 53.520 46.100 53.870 ;
        RECT 45.775 47.160 46.075 53.520 ;
        RECT 46.525 50.865 46.825 51.360 ;
        RECT 46.500 50.515 46.850 50.865 ;
        RECT 46.525 50.020 46.825 50.515 ;
        RECT 45.750 46.810 46.100 47.160 ;
        RECT 45.775 40.450 46.075 46.810 ;
        RECT 46.525 44.155 46.825 44.650 ;
        RECT 46.500 43.805 46.850 44.155 ;
        RECT 46.525 43.310 46.825 43.805 ;
        RECT 45.750 40.100 46.100 40.450 ;
        RECT 45.775 34.470 46.075 40.100 ;
        RECT 47.155 40.000 47.455 67.420 ;
        RECT 47.760 63.935 48.110 64.285 ;
        RECT 47.785 40.630 48.085 63.935 ;
        RECT 49.020 60.710 49.370 61.060 ;
        RECT 48.390 57.225 48.740 57.575 ;
        RECT 48.415 41.375 48.715 57.225 ;
        RECT 49.045 42.120 49.345 60.710 ;
        RECT 50.280 54.000 50.630 54.350 ;
        RECT 49.650 50.515 50.000 50.865 ;
        RECT 49.675 42.750 49.975 50.515 ;
        RECT 50.305 43.380 50.605 54.000 ;
        RECT 50.935 44.010 51.235 70.645 ;
        RECT 51.565 44.640 51.865 74.130 ;
        RECT 65.485 53.955 66.515 55.045 ;
        RECT 63.025 53.130 63.375 53.155 ;
        RECT 63.025 52.830 67.390 53.130 ;
        RECT 63.025 52.805 63.375 52.830 ;
        RECT 61.365 52.505 61.715 52.530 ;
        RECT 61.365 52.205 66.010 52.505 ;
        RECT 61.365 52.180 61.715 52.205 ;
        RECT 59.705 51.880 60.055 51.905 ;
        RECT 59.705 51.580 64.630 51.880 ;
        RECT 59.705 51.555 60.055 51.580 ;
        RECT 58.045 51.255 58.395 51.280 ;
        RECT 58.045 50.955 63.250 51.255 ;
        RECT 58.045 50.930 58.395 50.955 ;
        RECT 56.385 50.630 56.735 50.655 ;
        RECT 56.385 50.330 61.870 50.630 ;
        RECT 56.385 50.305 56.735 50.330 ;
        RECT 54.725 50.005 55.075 50.030 ;
        RECT 54.725 49.705 60.490 50.005 ;
        RECT 54.725 49.680 55.075 49.705 ;
        RECT 53.065 49.380 53.415 49.405 ;
        RECT 53.065 49.080 59.110 49.380 ;
        RECT 53.065 49.055 53.415 49.080 ;
        RECT 53.695 48.755 54.045 48.780 ;
        RECT 53.695 48.455 57.730 48.755 ;
        RECT 53.695 48.430 54.045 48.455 ;
        RECT 53.065 48.130 53.415 48.155 ;
        RECT 53.065 47.940 56.350 48.130 ;
        RECT 57.430 47.940 57.730 48.455 ;
        RECT 58.810 47.940 59.110 49.080 ;
        RECT 60.190 47.940 60.490 49.705 ;
        RECT 61.570 47.940 61.870 50.330 ;
        RECT 62.950 47.940 63.250 50.955 ;
        RECT 64.330 47.940 64.630 51.580 ;
        RECT 65.710 47.940 66.010 52.205 ;
        RECT 67.090 47.945 67.390 52.830 ;
        RECT 53.065 47.830 56.740 47.940 ;
        RECT 53.065 47.805 53.415 47.830 ;
        RECT 56.050 47.250 56.740 47.830 ;
        RECT 57.430 47.250 58.120 47.940 ;
        RECT 58.810 47.250 59.500 47.940 ;
        RECT 60.190 47.250 60.880 47.940 ;
        RECT 61.570 47.250 62.260 47.940 ;
        RECT 62.950 47.250 63.640 47.940 ;
        RECT 64.330 47.250 65.020 47.940 ;
        RECT 65.710 47.250 66.400 47.940 ;
        RECT 67.090 47.255 67.780 47.945 ;
        RECT 69.160 45.660 69.850 92.005 ;
        RECT 70.485 86.050 71.515 87.140 ;
        RECT 53.765 45.470 54.115 45.495 ;
        RECT 56.920 45.470 69.850 45.660 ;
        RECT 53.765 45.170 69.850 45.470 ;
        RECT 53.765 45.145 54.115 45.170 ;
        RECT 56.920 44.970 69.850 45.170 ;
        RECT 56.920 44.965 57.220 44.970 ;
        RECT 58.300 44.965 58.600 44.970 ;
        RECT 59.680 44.965 59.980 44.970 ;
        RECT 61.060 44.965 61.360 44.970 ;
        RECT 62.440 44.965 62.740 44.970 ;
        RECT 63.820 44.965 64.120 44.970 ;
        RECT 65.200 44.965 65.500 44.970 ;
        RECT 66.580 44.965 66.880 44.970 ;
        RECT 51.565 44.340 64.825 44.640 ;
        RECT 50.935 43.710 63.445 44.010 ;
        RECT 50.305 43.080 62.065 43.380 ;
        RECT 49.675 42.450 60.685 42.750 ;
        RECT 49.045 41.820 59.305 42.120 ;
        RECT 59.005 41.520 59.305 41.820 ;
        RECT 60.385 41.520 60.685 42.450 ;
        RECT 61.765 41.520 62.065 43.080 ;
        RECT 63.145 41.520 63.445 43.710 ;
        RECT 64.525 41.520 64.825 44.340 ;
        RECT 67.090 41.820 67.780 42.510 ;
        RECT 57.480 41.375 58.070 41.520 ;
        RECT 48.415 41.075 58.070 41.375 ;
        RECT 57.480 40.930 58.070 41.075 ;
        RECT 58.860 40.930 59.450 41.520 ;
        RECT 60.240 40.930 60.830 41.520 ;
        RECT 61.620 40.930 62.210 41.520 ;
        RECT 63.000 40.930 63.590 41.520 ;
        RECT 64.380 40.930 64.970 41.520 ;
        RECT 65.760 40.930 66.350 41.520 ;
        RECT 67.140 40.930 67.730 41.520 ;
        RECT 65.905 40.630 66.205 40.930 ;
        RECT 47.785 40.330 66.205 40.630 ;
        RECT 67.285 40.000 67.585 40.930 ;
        RECT 47.155 39.700 67.585 40.000 ;
        RECT 68.440 39.905 69.180 39.930 ;
        RECT 70.485 39.905 71.515 40.105 ;
        RECT 68.440 39.215 71.515 39.905 ;
        RECT 68.440 39.190 69.180 39.215 ;
        RECT 70.485 39.015 71.515 39.215 ;
        RECT 46.525 37.445 46.825 37.940 ;
        RECT 46.500 37.095 46.850 37.445 ;
        RECT 46.525 36.600 46.825 37.095 ;
        RECT 44.250 34.440 44.600 34.470 ;
        RECT 35.275 33.270 35.575 34.440 ;
        RECT 38.275 33.270 38.575 34.440 ;
        RECT 41.275 33.270 41.575 34.440 ;
        RECT 44.285 33.300 44.585 34.440 ;
        RECT 60.690 33.595 61.690 37.675 ;
        RECT 62.750 33.595 63.750 37.685 ;
        RECT 64.640 33.625 65.640 37.685 ;
        RECT 106.575 33.625 107.575 37.685 ;
        RECT 108.465 33.625 109.465 37.685 ;
        RECT 64.640 33.595 67.000 33.625 ;
        RECT 106.575 33.595 109.465 33.625 ;
        RECT 110.525 33.595 111.525 37.675 ;
        RECT 55.640 33.440 116.575 33.595 ;
        RECT 44.000 33.270 46.000 33.300 ;
        RECT 35.275 32.270 46.000 33.270 ;
        RECT 51.960 32.750 116.575 33.440 ;
        RECT 55.640 32.595 116.575 32.750 ;
        RECT 65.000 32.565 67.000 32.595 ;
        RECT 44.000 32.240 46.000 32.270 ;
        RECT 86.615 31.250 87.615 32.595 ;
        RECT 107.000 32.565 109.000 32.595 ;
        RECT 68.990 26.915 69.990 27.915 ;
        RECT 102.225 26.915 103.225 27.915 ;
        RECT 70.000 25.345 72.000 25.375 ;
        RECT 112.000 25.345 114.000 25.375 ;
        RECT 55.640 25.190 116.575 25.345 ;
        RECT 50.580 24.500 116.575 25.190 ;
        RECT 55.640 24.345 116.575 24.500 ;
        RECT 56.930 23.035 57.930 24.345 ;
        RECT 56.770 22.275 58.090 23.035 ;
        RECT 62.970 23.015 63.970 24.345 ;
        RECT 64.850 23.015 65.850 24.345 ;
        RECT 56.930 22.155 57.930 22.275 ;
        RECT 62.810 22.255 64.130 23.015 ;
        RECT 64.690 22.255 66.010 23.015 ;
        RECT 66.730 23.005 67.730 24.345 ;
        RECT 70.000 24.315 72.000 24.345 ;
        RECT 62.970 22.135 63.970 22.255 ;
        RECT 64.850 22.135 65.850 22.255 ;
        RECT 66.570 22.245 67.890 23.005 ;
        RECT 66.730 22.125 67.730 22.245 ;
        RECT 68.990 21.775 69.990 22.775 ;
        RECT 86.615 22.130 87.615 24.345 ;
        RECT 104.485 23.005 105.485 24.345 ;
        RECT 106.365 23.015 107.365 24.345 ;
        RECT 108.245 23.015 109.245 24.345 ;
        RECT 112.000 24.315 113.985 24.345 ;
        RECT 114.285 23.035 115.285 24.345 ;
        RECT 102.225 21.775 103.225 22.775 ;
        RECT 104.325 22.245 105.645 23.005 ;
        RECT 106.205 22.255 107.525 23.015 ;
        RECT 108.085 22.255 109.405 23.015 ;
        RECT 114.125 22.275 115.445 23.035 ;
        RECT 104.485 22.125 105.485 22.245 ;
        RECT 106.365 22.135 107.365 22.255 ;
        RECT 108.245 22.135 109.245 22.255 ;
        RECT 114.285 22.155 115.285 22.275 ;
        RECT 39.570 0.995 40.470 1.000 ;
        RECT 58.890 0.995 59.790 1.000 ;
        RECT 78.210 0.995 79.110 1.000 ;
        RECT 97.530 0.995 98.430 1.000 ;
        RECT 116.850 0.995 117.750 1.000 ;
        RECT 136.170 0.995 137.070 1.000 ;
        RECT 39.545 0.105 40.495 0.995 ;
        RECT 58.865 0.105 59.815 0.995 ;
        RECT 78.185 0.105 79.135 0.995 ;
        RECT 97.505 0.105 98.455 0.995 ;
        RECT 116.825 0.105 117.775 0.995 ;
        RECT 136.145 0.105 137.095 0.995 ;
        RECT 39.570 0.100 40.470 0.105 ;
        RECT 58.890 0.100 59.790 0.105 ;
        RECT 78.210 0.100 79.110 0.105 ;
        RECT 97.530 0.100 98.430 0.105 ;
        RECT 116.850 0.100 117.750 0.105 ;
        RECT 136.170 0.100 137.070 0.105 ;
      LAYER met4 ;
        RECT 20.535 225.085 20.550 225.090 ;
        RECT 15.005 224.760 15.030 225.085 ;
        RECT 15.330 224.760 15.355 225.085 ;
        RECT 15.005 224.735 15.355 224.760 ;
        RECT 17.765 224.760 17.790 225.085 ;
        RECT 18.090 224.760 18.115 225.085 ;
        RECT 17.765 224.735 18.115 224.760 ;
        RECT 20.525 224.760 20.550 225.085 ;
        RECT 20.850 225.085 20.865 225.090 ;
        RECT 20.850 224.760 20.875 225.085 ;
        RECT 20.525 224.735 20.875 224.760 ;
        RECT 23.285 224.760 23.310 225.085 ;
        RECT 23.610 224.760 23.635 225.085 ;
        RECT 23.285 224.735 23.635 224.760 ;
        RECT 26.045 224.760 26.070 225.085 ;
        RECT 26.370 224.760 26.395 225.085 ;
        RECT 26.045 224.735 26.395 224.760 ;
        RECT 28.805 224.760 28.830 225.085 ;
        RECT 29.130 224.760 29.155 225.085 ;
        RECT 28.805 224.735 29.155 224.760 ;
        RECT 31.565 224.760 31.590 225.085 ;
        RECT 31.890 224.760 31.915 225.085 ;
        RECT 31.565 224.735 31.915 224.760 ;
        RECT 34.325 224.760 34.350 225.085 ;
        RECT 34.650 224.760 34.675 225.085 ;
        RECT 34.325 224.735 34.675 224.760 ;
        RECT 37.085 224.760 37.110 225.085 ;
        RECT 37.410 224.760 37.435 225.085 ;
        RECT 37.085 224.735 37.435 224.760 ;
        RECT 39.845 224.760 39.870 225.085 ;
        RECT 40.170 224.760 40.195 225.085 ;
        RECT 39.845 224.735 40.195 224.760 ;
        RECT 42.605 224.760 42.630 225.085 ;
        RECT 42.930 224.760 42.955 225.085 ;
        RECT 42.605 224.735 42.955 224.760 ;
        RECT 45.365 224.760 45.390 225.085 ;
        RECT 45.690 224.760 45.715 225.085 ;
        RECT 45.365 224.735 45.715 224.760 ;
        RECT 48.125 224.760 48.150 225.085 ;
        RECT 48.450 224.760 48.475 225.085 ;
        RECT 48.125 224.735 48.475 224.760 ;
        RECT 50.885 224.760 50.910 225.085 ;
        RECT 51.210 224.760 51.235 225.085 ;
        RECT 50.885 224.735 51.235 224.760 ;
        RECT 53.645 224.760 53.670 225.085 ;
        RECT 53.970 224.760 53.995 225.085 ;
        RECT 53.645 224.735 53.995 224.760 ;
        RECT 56.405 224.760 56.430 225.085 ;
        RECT 56.730 224.760 56.755 225.085 ;
        RECT 56.405 224.735 56.755 224.760 ;
        RECT 59.165 224.760 59.190 225.085 ;
        RECT 59.490 224.760 59.515 225.085 ;
        RECT 59.165 224.735 59.515 224.760 ;
        RECT 61.925 224.760 61.950 225.085 ;
        RECT 62.250 224.760 62.275 225.085 ;
        RECT 61.925 224.735 62.275 224.760 ;
        RECT 64.685 224.760 64.710 225.085 ;
        RECT 65.010 224.760 65.035 225.085 ;
        RECT 64.685 224.735 65.035 224.760 ;
        RECT 67.445 224.760 67.470 225.085 ;
        RECT 67.770 224.760 67.795 225.085 ;
        RECT 67.445 224.735 67.795 224.760 ;
        RECT 70.205 224.760 70.230 225.085 ;
        RECT 70.530 224.760 70.555 225.085 ;
        RECT 70.205 224.735 70.555 224.760 ;
        RECT 72.965 224.760 72.990 225.085 ;
        RECT 73.290 224.760 73.315 225.085 ;
        RECT 72.965 224.735 73.315 224.760 ;
        RECT 75.725 224.760 75.750 225.085 ;
        RECT 76.050 224.760 76.075 225.085 ;
        RECT 75.725 224.735 76.075 224.760 ;
        RECT 78.485 224.760 78.510 225.085 ;
        RECT 78.810 224.760 78.835 225.085 ;
        RECT 98.130 224.760 98.155 225.085 ;
        RECT 103.325 224.760 103.350 225.085 ;
        RECT 103.650 224.760 103.675 225.085 ;
        RECT 78.485 224.735 78.835 224.760 ;
        RECT 103.325 224.735 103.675 224.760 ;
        RECT 106.085 224.760 106.110 225.085 ;
        RECT 106.410 224.760 106.435 225.085 ;
        RECT 106.085 224.735 106.435 224.760 ;
        RECT 108.845 224.760 108.870 225.085 ;
        RECT 109.170 224.760 109.195 225.085 ;
        RECT 108.845 224.735 109.195 224.760 ;
        RECT 111.605 224.760 111.630 225.085 ;
        RECT 111.930 224.760 111.955 225.085 ;
        RECT 111.605 224.735 111.955 224.760 ;
        RECT 114.365 224.760 114.390 225.085 ;
        RECT 114.690 224.760 114.715 225.085 ;
        RECT 114.365 224.735 114.715 224.760 ;
        RECT 117.125 224.760 117.150 225.085 ;
        RECT 117.450 224.760 117.475 225.085 ;
        RECT 117.125 224.735 117.475 224.760 ;
        RECT 119.885 224.760 119.910 225.085 ;
        RECT 120.210 224.760 120.235 225.085 ;
        RECT 119.885 224.735 120.235 224.760 ;
        RECT 122.645 224.760 122.670 225.085 ;
        RECT 122.970 224.760 122.995 225.085 ;
        RECT 122.645 224.735 122.995 224.760 ;
        RECT 38.995 207.805 39.000 208.165 ;
        RECT 41.000 207.805 41.005 208.165 ;
        RECT 43.995 207.805 44.000 208.165 ;
        RECT 46.000 207.805 46.005 208.165 ;
        RECT 48.995 207.805 49.000 208.165 ;
        RECT 51.000 207.805 51.005 208.165 ;
        RECT 64.995 207.805 65.000 208.165 ;
        RECT 67.000 207.805 67.005 208.165 ;
        RECT 69.995 207.805 70.000 208.165 ;
        RECT 72.000 207.805 72.005 208.165 ;
        RECT 74.995 207.805 75.000 208.165 ;
        RECT 77.000 207.805 77.005 208.165 ;
        RECT 20.995 206.380 21.000 206.740 ;
        RECT 23.000 206.380 23.005 206.740 ;
        RECT 106.995 206.300 107.000 206.660 ;
        RECT 109.000 206.300 109.005 206.660 ;
        RECT 111.995 206.300 112.000 206.660 ;
        RECT 114.000 206.300 114.005 206.660 ;
        RECT 116.995 206.300 117.000 206.660 ;
        RECT 119.000 206.300 119.005 206.660 ;
        RECT 38.995 202.145 39.000 202.505 ;
        RECT 41.000 202.145 41.005 202.505 ;
        RECT 43.995 202.145 44.000 202.505 ;
        RECT 46.000 202.145 46.005 202.505 ;
        RECT 48.995 202.145 49.000 202.505 ;
        RECT 51.000 202.145 51.005 202.505 ;
        RECT 64.995 202.145 65.000 202.505 ;
        RECT 67.000 202.145 67.005 202.505 ;
        RECT 69.995 202.145 70.000 202.505 ;
        RECT 72.000 202.145 72.005 202.505 ;
        RECT 74.995 202.145 75.000 202.505 ;
        RECT 77.000 202.145 77.005 202.505 ;
        RECT 38.995 201.095 39.000 201.455 ;
        RECT 41.000 201.095 41.005 201.455 ;
        RECT 43.995 201.095 44.000 201.455 ;
        RECT 46.000 201.095 46.005 201.455 ;
        RECT 48.995 201.095 49.000 201.455 ;
        RECT 51.000 201.095 51.005 201.455 ;
        RECT 64.995 201.095 65.000 201.455 ;
        RECT 67.000 201.095 67.005 201.455 ;
        RECT 69.995 201.095 70.000 201.455 ;
        RECT 72.000 201.095 72.005 201.455 ;
        RECT 74.995 201.095 75.000 201.455 ;
        RECT 77.000 201.095 77.005 201.455 ;
        RECT 15.995 200.715 16.000 201.075 ;
        RECT 18.000 200.715 18.015 201.075 ;
        RECT 106.995 200.640 107.000 201.000 ;
        RECT 109.000 200.640 109.005 201.000 ;
        RECT 111.995 200.640 112.000 201.000 ;
        RECT 114.000 200.640 114.005 201.000 ;
        RECT 116.995 200.640 117.000 201.000 ;
        RECT 119.000 200.640 119.005 201.000 ;
        RECT 38.995 195.435 39.000 195.795 ;
        RECT 41.000 195.435 41.005 195.795 ;
        RECT 43.995 195.435 44.000 195.795 ;
        RECT 46.000 195.435 46.005 195.795 ;
        RECT 48.995 195.435 49.000 195.795 ;
        RECT 51.000 195.435 51.005 195.795 ;
        RECT 64.995 195.435 65.000 195.795 ;
        RECT 67.000 195.435 67.005 195.795 ;
        RECT 69.995 195.435 70.000 195.795 ;
        RECT 72.000 195.435 72.005 195.795 ;
        RECT 74.995 195.435 75.000 195.795 ;
        RECT 77.000 195.435 77.005 195.795 ;
        RECT 106.995 188.835 107.000 189.195 ;
        RECT 109.000 188.835 109.005 189.195 ;
        RECT 111.995 188.835 112.000 189.195 ;
        RECT 114.000 188.835 114.005 189.195 ;
        RECT 116.995 188.835 117.000 189.195 ;
        RECT 119.000 188.835 119.005 189.195 ;
        RECT 38.995 183.630 39.000 183.990 ;
        RECT 41.000 183.630 41.005 183.990 ;
        RECT 43.995 183.630 44.000 183.990 ;
        RECT 46.000 183.630 46.005 183.990 ;
        RECT 48.995 183.630 49.000 183.990 ;
        RECT 51.000 183.630 51.005 183.990 ;
        RECT 64.995 183.630 65.000 183.990 ;
        RECT 67.000 183.630 67.005 183.990 ;
        RECT 69.995 183.630 70.000 183.990 ;
        RECT 72.000 183.630 72.005 183.990 ;
        RECT 74.995 183.630 75.000 183.990 ;
        RECT 77.000 183.630 77.005 183.990 ;
        RECT 106.995 183.175 107.000 183.535 ;
        RECT 109.000 183.175 109.005 183.535 ;
        RECT 111.995 183.175 112.000 183.535 ;
        RECT 114.000 183.175 114.005 183.535 ;
        RECT 116.995 183.175 117.000 183.535 ;
        RECT 119.000 183.175 119.005 183.535 ;
        RECT 106.995 182.125 107.000 182.485 ;
        RECT 109.000 182.125 109.005 182.485 ;
        RECT 111.995 182.125 112.000 182.485 ;
        RECT 114.000 182.125 114.005 182.485 ;
        RECT 116.995 182.125 117.000 182.485 ;
        RECT 119.000 182.125 119.005 182.485 ;
        RECT 38.995 177.970 39.000 178.330 ;
        RECT 41.000 177.970 41.005 178.330 ;
        RECT 43.995 177.970 44.000 178.330 ;
        RECT 46.000 177.970 46.005 178.330 ;
        RECT 48.995 177.970 49.000 178.330 ;
        RECT 51.000 177.970 51.005 178.330 ;
        RECT 64.995 177.970 65.000 178.330 ;
        RECT 67.000 177.970 67.005 178.330 ;
        RECT 69.995 177.970 70.000 178.330 ;
        RECT 72.000 177.970 72.005 178.330 ;
        RECT 74.995 177.970 75.000 178.330 ;
        RECT 77.000 177.970 77.005 178.330 ;
        RECT 38.995 176.920 39.000 177.280 ;
        RECT 41.000 176.920 41.005 177.280 ;
        RECT 43.995 176.920 44.000 177.280 ;
        RECT 46.000 176.920 46.005 177.280 ;
        RECT 48.995 176.920 49.000 177.280 ;
        RECT 51.000 176.920 51.005 177.280 ;
        RECT 106.995 176.465 107.000 176.825 ;
        RECT 109.000 176.465 109.005 176.825 ;
        RECT 111.995 176.465 112.000 176.825 ;
        RECT 114.000 176.465 114.005 176.825 ;
        RECT 116.995 176.465 117.000 176.825 ;
        RECT 119.000 176.465 119.005 176.825 ;
        RECT 38.995 145.690 39.000 146.050 ;
        RECT 41.000 145.690 41.005 146.050 ;
        RECT 43.995 145.690 44.000 146.050 ;
        RECT 46.000 145.690 46.005 146.050 ;
        RECT 48.995 145.690 49.000 146.050 ;
        RECT 51.000 145.690 51.005 146.050 ;
        RECT 64.995 145.690 65.000 146.050 ;
        RECT 67.000 145.690 67.005 146.050 ;
        RECT 69.995 145.690 70.000 146.050 ;
        RECT 72.000 145.690 72.005 146.050 ;
        RECT 74.995 145.690 75.000 146.050 ;
        RECT 77.000 145.690 77.005 146.050 ;
        RECT 38.995 144.190 39.000 144.550 ;
        RECT 41.000 144.190 41.005 144.550 ;
        RECT 43.995 144.190 44.000 144.550 ;
        RECT 46.000 144.190 46.005 144.550 ;
        RECT 48.995 144.190 49.000 144.550 ;
        RECT 51.000 144.190 51.005 144.550 ;
        RECT 64.995 144.190 65.000 144.550 ;
        RECT 67.000 144.190 67.005 144.550 ;
        RECT 69.995 144.190 70.000 144.550 ;
        RECT 72.000 144.190 72.005 144.550 ;
        RECT 74.995 144.190 75.000 144.550 ;
        RECT 77.000 144.190 77.005 144.550 ;
        RECT 38.995 142.690 39.000 143.050 ;
        RECT 41.000 142.690 41.005 143.050 ;
        RECT 43.995 142.690 44.000 143.050 ;
        RECT 46.000 142.690 46.005 143.050 ;
        RECT 48.995 142.690 49.000 143.050 ;
        RECT 51.000 142.690 51.005 143.050 ;
        RECT 64.995 142.690 65.000 143.050 ;
        RECT 67.000 142.690 67.005 143.050 ;
        RECT 69.995 142.690 70.000 143.050 ;
        RECT 72.000 142.690 72.005 143.050 ;
        RECT 74.995 142.690 75.000 143.050 ;
        RECT 77.000 142.690 77.005 143.050 ;
        RECT 38.995 141.190 39.000 141.550 ;
        RECT 41.000 141.190 41.005 141.550 ;
        RECT 43.995 141.190 44.000 141.550 ;
        RECT 46.000 141.190 46.005 141.550 ;
        RECT 48.995 141.190 49.000 141.550 ;
        RECT 51.000 141.190 51.005 141.550 ;
        RECT 64.995 141.190 65.000 141.550 ;
        RECT 67.000 141.190 67.005 141.550 ;
        RECT 69.995 141.190 70.000 141.550 ;
        RECT 72.000 141.190 72.005 141.550 ;
        RECT 74.995 141.190 75.000 141.550 ;
        RECT 77.000 141.190 77.005 141.550 ;
        RECT 38.995 139.690 39.000 140.050 ;
        RECT 41.000 139.690 41.005 140.050 ;
        RECT 43.995 139.690 44.000 140.050 ;
        RECT 46.000 139.690 46.005 140.050 ;
        RECT 48.995 139.690 49.000 140.050 ;
        RECT 51.000 139.690 51.005 140.050 ;
        RECT 64.995 139.690 65.000 140.050 ;
        RECT 67.000 139.690 67.005 140.050 ;
        RECT 69.995 139.690 70.000 140.050 ;
        RECT 72.000 139.690 72.005 140.050 ;
        RECT 74.995 139.690 75.000 140.050 ;
        RECT 77.000 139.690 77.005 140.050 ;
        RECT 38.995 138.190 39.000 138.550 ;
        RECT 41.000 138.190 41.005 138.550 ;
        RECT 43.995 138.190 44.000 138.550 ;
        RECT 46.000 138.190 46.005 138.550 ;
        RECT 48.995 138.190 49.000 138.550 ;
        RECT 51.000 138.190 51.005 138.550 ;
        RECT 64.995 138.190 65.000 138.550 ;
        RECT 67.000 138.190 67.005 138.550 ;
        RECT 69.995 138.190 70.000 138.550 ;
        RECT 72.000 138.190 72.005 138.550 ;
        RECT 74.995 138.190 75.000 138.550 ;
        RECT 77.000 138.190 77.005 138.550 ;
        RECT 38.995 136.690 39.000 137.050 ;
        RECT 41.000 136.690 41.005 137.050 ;
        RECT 43.995 136.690 44.000 137.050 ;
        RECT 46.000 136.690 46.005 137.050 ;
        RECT 48.995 136.690 49.000 137.050 ;
        RECT 51.000 136.690 51.005 137.050 ;
        RECT 64.995 136.690 65.000 137.050 ;
        RECT 67.000 136.690 67.005 137.050 ;
        RECT 69.995 136.690 70.000 137.050 ;
        RECT 72.000 136.690 72.005 137.050 ;
        RECT 74.995 136.690 75.000 137.050 ;
        RECT 77.000 136.690 77.005 137.050 ;
        RECT 38.995 135.190 39.000 135.550 ;
        RECT 41.000 135.190 41.005 135.550 ;
        RECT 43.995 135.190 44.000 135.550 ;
        RECT 46.000 135.190 46.005 135.550 ;
        RECT 48.995 135.190 49.000 135.550 ;
        RECT 51.000 135.190 51.005 135.550 ;
        RECT 64.995 135.190 65.000 135.550 ;
        RECT 67.000 135.190 67.005 135.550 ;
        RECT 69.995 135.190 70.000 135.550 ;
        RECT 72.000 135.190 72.005 135.550 ;
        RECT 74.995 135.190 75.000 135.550 ;
        RECT 77.000 135.190 77.005 135.550 ;
        RECT 38.995 133.690 39.000 134.050 ;
        RECT 41.000 133.690 41.005 134.050 ;
        RECT 43.995 133.690 44.000 134.050 ;
        RECT 46.000 133.690 46.005 134.050 ;
        RECT 48.995 133.690 49.000 134.050 ;
        RECT 51.000 133.690 51.005 134.050 ;
        RECT 64.995 133.690 65.000 134.050 ;
        RECT 67.000 133.690 67.005 134.050 ;
        RECT 69.995 133.690 70.000 134.050 ;
        RECT 72.000 133.690 72.005 134.050 ;
        RECT 74.995 133.690 75.000 134.050 ;
        RECT 77.000 133.690 77.005 134.050 ;
        RECT 38.995 120.995 39.000 123.005 ;
        RECT 41.000 120.995 41.005 123.005 ;
        RECT 64.995 120.995 65.000 123.005 ;
        RECT 67.000 120.995 67.005 123.005 ;
        RECT 106.995 120.995 107.000 123.005 ;
        RECT 109.000 120.995 109.005 123.005 ;
        RECT 15.995 115.995 16.000 118.005 ;
        RECT 18.000 115.995 18.005 118.005 ;
        RECT 43.995 115.995 44.000 118.005 ;
        RECT 46.000 115.995 46.005 118.005 ;
        RECT 69.995 115.995 70.000 118.005 ;
        RECT 72.000 115.995 72.005 118.005 ;
        RECT 111.995 115.995 112.000 118.005 ;
        RECT 114.000 115.995 114.005 118.005 ;
        RECT 20.995 110.995 21.000 113.005 ;
        RECT 23.000 110.995 23.005 113.005 ;
        RECT 48.995 110.995 49.000 113.005 ;
        RECT 51.000 110.995 51.005 113.005 ;
        RECT 74.995 110.995 75.000 113.005 ;
        RECT 77.000 110.995 77.005 113.005 ;
        RECT 116.995 110.995 117.000 113.005 ;
        RECT 119.000 110.995 119.005 113.005 ;
        RECT 38.995 102.005 39.000 103.015 ;
        RECT 41.000 102.005 41.005 103.015 ;
        RECT 72.000 85.905 72.005 87.285 ;
        RECT 43.995 32.265 44.000 33.275 ;
        RECT 46.000 32.265 46.005 33.275 ;
        RECT 64.995 32.590 65.000 33.600 ;
        RECT 67.000 32.590 67.005 33.600 ;
        RECT 106.995 32.590 107.000 33.600 ;
        RECT 109.000 32.590 109.005 33.600 ;
        RECT 69.995 24.340 70.000 25.350 ;
        RECT 72.000 24.340 72.005 25.350 ;
        RECT 111.995 24.340 112.000 25.350 ;
        RECT 114.000 24.340 114.005 25.350 ;
  END
END tt_um_htfab_hybrid
END LIBRARY

