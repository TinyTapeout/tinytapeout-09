VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_snn_with_delays_paolaunisa
  CLASS BLOCK ;
  FOREIGN tt_um_snn_with_delays_paolaunisa ;
  ORIGIN 0.000 0.000 ;
  SIZE 1378.160 BY 225.760 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.580 2.480 23.180 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.450 2.480 62.050 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.320 2.480 100.920 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.190 2.480 139.790 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.060 2.480 178.660 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 215.930 2.480 217.530 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.800 2.480 256.400 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 293.670 2.480 295.270 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.540 2.480 334.140 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.410 2.480 373.010 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.280 2.480 411.880 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 449.150 2.480 450.750 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.020 2.480 489.620 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 526.890 2.480 528.490 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 565.760 2.480 567.360 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.630 2.480 606.230 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 643.500 2.480 645.100 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 682.370 2.480 683.970 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.240 2.480 722.840 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 760.110 2.480 761.710 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 798.980 2.480 800.580 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.850 2.480 839.450 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 876.720 2.480 878.320 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 915.590 2.480 917.190 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.460 2.480 956.060 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 993.330 2.480 994.930 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.200 2.480 1033.800 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.070 2.480 1072.670 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1109.940 2.480 1111.540 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1148.810 2.480 1150.410 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1187.680 2.480 1189.280 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1226.550 2.480 1228.150 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1265.420 2.480 1267.020 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.290 2.480 1305.890 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1343.160 2.480 1344.760 223.280 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.150 2.480 58.750 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.020 2.480 97.620 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.890 2.480 136.490 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 173.760 2.480 175.360 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 212.630 2.480 214.230 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.500 2.480 253.100 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.370 2.480 291.970 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 329.240 2.480 330.840 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.110 2.480 369.710 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.980 2.480 408.580 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 445.850 2.480 447.450 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.720 2.480 486.320 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.590 2.480 525.190 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 562.460 2.480 564.060 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.330 2.480 602.930 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 640.200 2.480 641.800 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 679.070 2.480 680.670 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 717.940 2.480 719.540 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 756.810 2.480 758.410 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 795.680 2.480 797.280 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 834.550 2.480 836.150 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 873.420 2.480 875.020 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 912.290 2.480 913.890 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.160 2.480 952.760 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 990.030 2.480 991.630 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1028.900 2.480 1030.500 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1067.770 2.480 1069.370 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1106.640 2.480 1108.240 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.510 2.480 1147.110 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.380 2.480 1185.980 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.250 2.480 1224.850 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1262.120 2.480 1263.720 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1300.990 2.480 1302.590 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1339.860 2.480 1341.460 223.280 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 2.635 1375.590 223.230 ;
      LAYER li1 ;
        RECT 2.760 2.635 1375.400 223.125 ;
      LAYER met1 ;
        RECT 2.760 0.040 1375.400 225.720 ;
      LAYER met2 ;
        RECT 11.140 0.010 1366.560 225.750 ;
      LAYER met3 ;
        RECT 14.325 0.175 1361.075 225.585 ;
      LAYER met4 ;
        RECT 24.215 224.360 30.270 225.585 ;
        RECT 31.370 224.360 33.030 225.585 ;
        RECT 34.130 224.360 35.790 225.585 ;
        RECT 36.890 224.360 38.550 225.585 ;
        RECT 39.650 224.360 41.310 225.585 ;
        RECT 42.410 224.360 44.070 225.585 ;
        RECT 45.170 224.360 46.830 225.585 ;
        RECT 47.930 224.360 49.590 225.585 ;
        RECT 50.690 224.360 52.350 225.585 ;
        RECT 53.450 224.360 55.110 225.585 ;
        RECT 56.210 224.360 57.870 225.585 ;
        RECT 58.970 224.360 60.630 225.585 ;
        RECT 61.730 224.360 63.390 225.585 ;
        RECT 64.490 224.360 66.150 225.585 ;
        RECT 67.250 224.360 68.910 225.585 ;
        RECT 70.010 224.360 71.670 225.585 ;
        RECT 72.770 224.360 74.430 225.585 ;
        RECT 75.530 224.360 77.190 225.585 ;
        RECT 78.290 224.360 79.950 225.585 ;
        RECT 81.050 224.360 82.710 225.585 ;
        RECT 83.810 224.360 85.470 225.585 ;
        RECT 86.570 224.360 88.230 225.585 ;
        RECT 89.330 224.360 90.990 225.585 ;
        RECT 92.090 224.360 93.750 225.585 ;
        RECT 94.850 224.360 96.510 225.585 ;
        RECT 97.610 224.360 99.270 225.585 ;
        RECT 100.370 224.360 102.030 225.585 ;
        RECT 103.130 224.360 104.790 225.585 ;
        RECT 105.890 224.360 107.550 225.585 ;
        RECT 108.650 224.360 110.310 225.585 ;
        RECT 111.410 224.360 113.070 225.585 ;
        RECT 114.170 224.360 115.830 225.585 ;
        RECT 116.930 224.360 118.590 225.585 ;
        RECT 119.690 224.360 121.350 225.585 ;
        RECT 122.450 224.360 124.110 225.585 ;
        RECT 125.210 224.360 126.870 225.585 ;
        RECT 127.970 224.360 129.630 225.585 ;
        RECT 130.730 224.360 132.390 225.585 ;
        RECT 133.490 224.360 135.150 225.585 ;
        RECT 136.250 224.360 137.910 225.585 ;
        RECT 139.010 224.360 140.670 225.585 ;
        RECT 141.770 224.360 143.430 225.585 ;
        RECT 144.530 224.360 146.190 225.585 ;
        RECT 147.290 224.360 1256.425 225.585 ;
        RECT 24.215 223.680 1256.425 224.360 ;
        RECT 24.215 2.080 56.750 223.680 ;
        RECT 59.150 2.080 60.050 223.680 ;
        RECT 62.450 2.080 95.620 223.680 ;
        RECT 98.020 2.080 98.920 223.680 ;
        RECT 101.320 2.080 134.490 223.680 ;
        RECT 136.890 2.080 137.790 223.680 ;
        RECT 140.190 2.080 173.360 223.680 ;
        RECT 175.760 2.080 176.660 223.680 ;
        RECT 179.060 2.080 212.230 223.680 ;
        RECT 214.630 2.080 215.530 223.680 ;
        RECT 217.930 2.080 251.100 223.680 ;
        RECT 253.500 2.080 254.400 223.680 ;
        RECT 256.800 2.080 289.970 223.680 ;
        RECT 292.370 2.080 293.270 223.680 ;
        RECT 295.670 2.080 328.840 223.680 ;
        RECT 331.240 2.080 332.140 223.680 ;
        RECT 334.540 2.080 367.710 223.680 ;
        RECT 370.110 2.080 371.010 223.680 ;
        RECT 373.410 2.080 406.580 223.680 ;
        RECT 408.980 2.080 409.880 223.680 ;
        RECT 412.280 2.080 445.450 223.680 ;
        RECT 447.850 2.080 448.750 223.680 ;
        RECT 451.150 2.080 484.320 223.680 ;
        RECT 486.720 2.080 487.620 223.680 ;
        RECT 490.020 2.080 523.190 223.680 ;
        RECT 525.590 2.080 526.490 223.680 ;
        RECT 528.890 2.080 562.060 223.680 ;
        RECT 564.460 2.080 565.360 223.680 ;
        RECT 567.760 2.080 600.930 223.680 ;
        RECT 603.330 2.080 604.230 223.680 ;
        RECT 606.630 2.080 639.800 223.680 ;
        RECT 642.200 2.080 643.100 223.680 ;
        RECT 645.500 2.080 678.670 223.680 ;
        RECT 681.070 2.080 681.970 223.680 ;
        RECT 684.370 2.080 717.540 223.680 ;
        RECT 719.940 2.080 720.840 223.680 ;
        RECT 723.240 2.080 756.410 223.680 ;
        RECT 758.810 2.080 759.710 223.680 ;
        RECT 762.110 2.080 795.280 223.680 ;
        RECT 797.680 2.080 798.580 223.680 ;
        RECT 800.980 2.080 834.150 223.680 ;
        RECT 836.550 2.080 837.450 223.680 ;
        RECT 839.850 2.080 873.020 223.680 ;
        RECT 875.420 2.080 876.320 223.680 ;
        RECT 878.720 2.080 911.890 223.680 ;
        RECT 914.290 2.080 915.190 223.680 ;
        RECT 917.590 2.080 950.760 223.680 ;
        RECT 953.160 2.080 954.060 223.680 ;
        RECT 956.460 2.080 989.630 223.680 ;
        RECT 992.030 2.080 992.930 223.680 ;
        RECT 995.330 2.080 1028.500 223.680 ;
        RECT 1030.900 2.080 1031.800 223.680 ;
        RECT 1034.200 2.080 1067.370 223.680 ;
        RECT 1069.770 2.080 1070.670 223.680 ;
        RECT 1073.070 2.080 1106.240 223.680 ;
        RECT 1108.640 2.080 1109.540 223.680 ;
        RECT 1111.940 2.080 1145.110 223.680 ;
        RECT 1147.510 2.080 1148.410 223.680 ;
        RECT 1150.810 2.080 1183.980 223.680 ;
        RECT 1186.380 2.080 1187.280 223.680 ;
        RECT 1189.680 2.080 1222.850 223.680 ;
        RECT 1225.250 2.080 1226.150 223.680 ;
        RECT 1228.550 2.080 1256.425 223.680 ;
        RECT 24.215 0.175 1256.425 2.080 ;
  END
END tt_um_snn_with_delays_paolaunisa
END LIBRARY

