VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_r2r_dac
  CLASS BLOCK ;
  FOREIGN tt_um_r2r_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 115.590 199.020 116.090 199.110 ;
        RECT 121.980 199.090 122.480 199.110 ;
        RECT 103.980 198.700 104.480 198.790 ;
        RECT 110.370 198.770 110.870 198.790 ;
        RECT 102.850 196.200 105.360 198.700 ;
        RECT 108.880 196.270 111.390 198.770 ;
        RECT 114.460 196.520 116.970 199.020 ;
        RECT 120.490 196.590 123.000 199.090 ;
        RECT 127.600 199.020 128.100 199.110 ;
        RECT 133.990 199.090 134.490 199.110 ;
        RECT 126.470 196.520 128.980 199.020 ;
        RECT 132.500 196.590 135.010 199.090 ;
        RECT 138.730 199.030 139.230 199.120 ;
        RECT 145.120 199.100 145.620 199.120 ;
        RECT 137.600 196.530 140.110 199.030 ;
        RECT 143.630 196.600 146.140 199.100 ;
        RECT 138.660 182.480 139.160 182.570 ;
        RECT 145.050 182.550 145.550 182.570 ;
        RECT 103.340 182.200 103.840 182.220 ;
        RECT 102.820 179.700 105.330 182.200 ;
        RECT 109.730 182.130 110.230 182.220 ;
        RECT 108.850 179.630 111.360 182.130 ;
        RECT 126.650 182.080 127.150 182.170 ;
        RECT 133.040 182.150 133.540 182.170 ;
        RECT 115.650 181.890 116.150 181.980 ;
        RECT 122.040 181.960 122.540 181.980 ;
        RECT 114.520 179.390 117.030 181.890 ;
        RECT 120.550 179.460 123.060 181.960 ;
        RECT 125.520 179.580 128.030 182.080 ;
        RECT 131.550 179.650 134.060 182.150 ;
        RECT 137.530 179.980 140.040 182.480 ;
        RECT 143.560 180.050 146.070 182.550 ;
        RECT 91.970 164.630 92.470 164.650 ;
        RECT 91.450 162.130 93.960 164.630 ;
        RECT 98.360 164.560 98.860 164.650 ;
        RECT 103.080 164.620 103.580 164.640 ;
        RECT 97.480 162.060 99.990 164.560 ;
        RECT 102.560 162.120 105.070 164.620 ;
        RECT 109.470 164.550 109.970 164.640 ;
        RECT 114.110 164.560 114.610 164.580 ;
        RECT 108.590 162.050 111.100 164.550 ;
        RECT 113.590 162.060 116.100 164.560 ;
        RECT 120.500 164.490 121.000 164.580 ;
        RECT 124.590 164.510 125.090 164.530 ;
        RECT 119.620 161.990 122.130 164.490 ;
        RECT 124.070 162.010 126.580 164.510 ;
        RECT 130.980 164.440 131.480 164.530 ;
        RECT 134.660 164.520 135.160 164.540 ;
        RECT 130.100 161.940 132.610 164.440 ;
        RECT 134.140 162.020 136.650 164.520 ;
        RECT 141.050 164.450 141.550 164.540 ;
        RECT 140.170 161.950 142.680 164.450 ;
      LAYER met1 ;
        RECT 131.740 218.100 133.060 218.150 ;
        RECT 129.450 217.000 130.850 218.100 ;
        RECT 131.740 217.460 133.390 218.100 ;
        RECT 131.740 217.280 133.580 217.460 ;
        RECT 129.260 216.670 130.960 217.000 ;
        RECT 131.630 216.950 133.580 217.280 ;
        RECT 99.900 215.650 130.960 216.670 ;
        RECT 99.900 197.870 100.920 215.650 ;
        RECT 129.260 215.600 130.960 215.650 ;
        RECT 131.740 216.490 133.580 216.950 ;
        RECT 135.150 216.740 136.550 218.050 ;
        RECT 138.040 217.700 139.440 218.110 ;
        RECT 137.950 216.960 139.620 217.700 ;
        RECT 138.000 216.760 139.420 216.960 ;
        RECT 131.740 214.310 133.060 216.490 ;
        RECT 112.510 212.990 133.060 214.310 ;
        RECT 102.430 197.870 105.820 198.960 ;
        RECT 99.900 196.850 105.820 197.870 ;
        RECT 102.430 195.880 105.820 196.850 ;
        RECT 108.770 196.390 111.460 198.850 ;
        RECT 112.510 198.300 113.830 212.990 ;
        RECT 135.310 212.740 136.450 216.740 ;
        RECT 138.250 216.500 138.950 216.760 ;
        RECT 124.990 211.600 136.450 212.740 ;
        RECT 138.340 212.040 138.800 216.500 ;
        RECT 114.250 198.300 117.130 199.170 ;
        RECT 112.510 196.980 117.130 198.300 ;
        RECT 108.740 195.490 111.500 196.390 ;
        RECT 114.250 196.380 117.130 196.980 ;
        RECT 120.380 196.540 123.070 199.170 ;
        RECT 124.990 198.480 126.130 211.600 ;
        RECT 137.240 211.580 138.800 212.040 ;
        RECT 126.300 198.480 129.070 199.140 ;
        RECT 124.990 197.340 129.070 198.480 ;
        RECT 120.470 195.970 123.010 196.540 ;
        RECT 126.300 196.410 129.070 197.340 ;
        RECT 132.390 197.190 135.080 199.170 ;
        RECT 132.360 196.020 135.080 197.190 ;
        RECT 137.250 199.150 137.695 211.580 ;
        RECT 137.250 196.760 140.210 199.150 ;
        RECT 137.450 196.470 140.210 196.760 ;
        RECT 143.520 196.580 146.210 199.180 ;
        RECT 100.700 195.010 111.500 195.490 ;
        RECT 100.670 194.420 111.500 195.010 ;
        RECT 113.350 194.990 123.010 195.970 ;
        RECT 124.370 195.020 135.080 196.020 ;
        RECT 143.510 196.010 146.330 196.580 ;
        RECT 136.420 195.020 146.370 196.010 ;
        RECT 100.670 194.410 111.460 194.420 ;
        RECT 100.670 182.280 102.780 194.410 ;
        RECT 100.670 181.700 105.440 182.280 ;
        RECT 100.640 180.440 105.440 181.700 ;
        RECT 102.750 179.650 105.440 180.440 ;
        RECT 108.780 179.920 111.470 182.210 ;
        RECT 113.390 181.970 115.430 194.990 ;
        RECT 120.470 194.940 123.010 194.990 ;
        RECT 124.390 194.810 126.660 195.020 ;
        RECT 136.400 194.990 146.370 195.020 ;
        RECT 124.390 182.160 126.420 194.810 ;
        RECT 136.400 182.560 138.390 194.990 ;
        RECT 113.390 180.950 117.100 181.970 ;
        RECT 108.720 178.490 113.180 179.920 ;
        RECT 114.410 179.340 117.100 180.950 ;
        RECT 120.440 180.520 123.130 182.040 ;
        RECT 124.390 180.980 128.100 182.160 ;
        RECT 90.780 161.710 94.500 164.890 ;
        RECT 97.410 164.110 100.100 164.640 ;
        RECT 102.490 164.110 105.180 164.700 ;
        RECT 97.410 162.450 105.180 164.110 ;
        RECT 97.410 162.010 100.100 162.450 ;
        RECT 102.490 162.070 105.180 162.450 ;
        RECT 108.520 163.900 111.210 164.630 ;
        RECT 111.660 163.900 113.030 178.490 ;
        RECT 115.140 164.640 116.930 179.340 ;
        RECT 120.370 179.070 123.950 180.520 ;
        RECT 125.410 179.530 128.100 180.980 ;
        RECT 131.440 179.600 134.130 182.230 ;
        RECT 136.400 180.020 140.110 182.560 ;
        RECT 143.450 180.020 146.140 182.630 ;
        RECT 137.420 179.930 140.110 180.020 ;
        RECT 143.420 180.000 146.140 180.020 ;
        RECT 132.550 179.150 134.380 179.600 ;
        RECT 120.370 178.950 123.970 179.070 ;
        RECT 122.180 164.800 123.970 178.950 ;
        RECT 113.520 164.430 116.930 164.640 ;
        RECT 121.890 164.590 124.120 164.800 ;
        RECT 132.590 164.600 134.380 179.150 ;
        RECT 143.420 164.720 146.110 180.000 ;
        RECT 121.890 164.570 126.690 164.590 ;
        RECT 113.520 163.900 116.210 164.430 ;
        RECT 108.520 162.520 116.210 163.900 ;
        RECT 108.520 162.000 111.210 162.520 ;
        RECT 113.520 162.010 116.210 162.520 ;
        RECT 119.550 162.420 126.690 164.570 ;
        RECT 132.590 164.520 136.760 164.600 ;
        RECT 119.550 161.940 122.240 162.420 ;
        RECT 124.000 161.960 126.690 162.420 ;
        RECT 130.030 162.430 136.760 164.520 ;
        RECT 130.030 161.890 132.720 162.430 ;
        RECT 134.070 161.970 136.760 162.430 ;
        RECT 139.610 163.705 146.110 164.720 ;
        RECT 139.610 161.995 151.245 163.705 ;
        RECT 91.525 159.860 93.875 161.710 ;
        RECT 139.610 161.160 146.110 161.995 ;
        RECT 139.610 161.150 143.590 161.160 ;
        RECT 91.525 157.510 110.380 159.860 ;
        RECT 108.030 157.210 110.380 157.510 ;
        RECT 105.530 153.060 112.480 157.210 ;
        RECT 149.535 155.770 151.245 161.995 ;
        RECT 147.800 154.650 152.830 155.770 ;
        RECT 147.310 151.110 153.770 154.650 ;
      LAYER met2 ;
        RECT 129.120 218.810 131.170 220.760 ;
        RECT 129.690 217.990 130.610 218.810 ;
        RECT 131.950 218.720 134.000 220.670 ;
        RECT 132.380 217.990 133.300 218.720 ;
        RECT 135.080 218.520 137.130 220.470 ;
        RECT 129.540 216.860 130.710 217.990 ;
        RECT 132.080 217.620 133.300 217.990 ;
        RECT 135.440 217.940 136.360 218.520 ;
        RECT 137.630 218.500 139.680 220.450 ;
        RECT 138.300 218.000 139.220 218.500 ;
        RECT 132.080 216.860 133.250 217.620 ;
        RECT 135.240 216.810 136.410 217.940 ;
        RECT 138.130 216.870 139.300 218.000 ;
        RECT 105.120 152.240 113.550 157.430 ;
        RECT 107.920 151.200 111.530 152.240 ;
        RECT 147.570 151.300 153.360 154.350 ;
        RECT 105.580 147.270 113.530 151.200 ;
        RECT 148.120 149.780 152.960 151.300 ;
        RECT 147.390 147.140 153.840 149.780 ;
      LAYER met3 ;
        RECT 135.000 224.750 136.210 224.760 ;
        RECT 129.600 223.840 130.600 224.750 ;
        RECT 129.970 220.660 130.330 223.840 ;
        RECT 132.350 223.540 133.500 224.750 ;
        RECT 134.900 223.550 136.260 224.750 ;
        RECT 137.750 224.000 139.060 224.750 ;
        RECT 137.750 223.800 139.050 224.000 ;
        RECT 129.170 218.860 130.970 220.660 ;
        RECT 132.780 220.570 133.140 223.540 ;
        RECT 132.000 218.770 133.800 220.570 ;
        RECT 135.245 220.370 135.695 223.550 ;
        RECT 135.130 218.570 136.930 220.370 ;
        RECT 138.150 220.350 138.470 223.800 ;
        RECT 137.680 218.550 139.480 220.350 ;
        RECT 105.120 146.850 114.200 151.420 ;
        RECT 107.470 144.360 111.120 146.850 ;
        RECT 147.010 146.190 154.370 149.980 ;
        RECT 148.300 144.860 153.170 146.190 ;
        RECT 105.820 142.050 113.240 144.360 ;
        RECT 147.160 141.790 154.320 144.860 ;
        RECT 147.570 141.130 154.310 141.790 ;
      LAYER met4 ;
        RECT 91.300 224.800 91.390 225.100 ;
        RECT 96.600 224.800 96.910 225.290 ;
        RECT 4.975 224.760 30.670 224.800 ;
        RECT 30.970 224.760 33.430 224.800 ;
        RECT 33.730 224.760 36.190 224.800 ;
        RECT 36.490 224.760 38.950 224.800 ;
        RECT 39.250 224.760 41.710 224.800 ;
        RECT 42.010 224.760 44.470 224.800 ;
        RECT 44.770 224.760 47.230 224.800 ;
        RECT 47.530 224.760 49.990 224.800 ;
        RECT 50.290 224.760 52.750 224.800 ;
        RECT 53.050 224.760 55.510 224.800 ;
        RECT 55.810 224.760 58.270 224.800 ;
        RECT 58.570 224.760 61.030 224.800 ;
        RECT 61.330 224.760 63.790 224.800 ;
        RECT 64.090 224.760 66.550 224.800 ;
        RECT 66.850 224.760 69.310 224.800 ;
        RECT 69.610 224.760 72.070 224.800 ;
        RECT 72.370 224.760 74.830 224.800 ;
        RECT 75.130 224.760 77.590 224.800 ;
        RECT 77.890 224.760 80.350 224.800 ;
        RECT 80.650 224.760 83.110 224.800 ;
        RECT 83.410 224.760 85.870 224.800 ;
        RECT 86.170 224.760 88.630 224.800 ;
        RECT 88.930 224.760 91.390 224.800 ;
        RECT 91.690 224.760 94.150 224.800 ;
        RECT 94.450 224.760 95.330 224.800 ;
        RECT 4.975 224.450 95.330 224.760 ;
        RECT 96.010 224.760 96.910 224.800 ;
        RECT 97.210 224.800 97.540 225.240 ;
        RECT 97.210 224.760 98.660 224.800 ;
        RECT 96.010 224.450 98.660 224.760 ;
        RECT 99.340 224.760 99.670 224.800 ;
        RECT 99.970 224.760 100.980 224.800 ;
        RECT 99.340 224.450 100.980 224.760 ;
        RECT 101.660 224.760 102.430 224.800 ;
        RECT 102.730 224.760 103.900 224.800 ;
        RECT 101.660 224.450 103.900 224.760 ;
        RECT 104.580 224.760 105.190 224.800 ;
        RECT 105.490 224.760 106.540 224.800 ;
        RECT 104.580 224.450 106.540 224.760 ;
        RECT 107.220 224.760 107.950 224.800 ;
        RECT 108.250 224.760 109.370 224.800 ;
        RECT 107.220 224.450 109.370 224.760 ;
        RECT 110.050 224.760 110.710 224.800 ;
        RECT 111.010 224.760 111.910 224.800 ;
        RECT 110.050 224.450 111.910 224.760 ;
        RECT 112.590 224.760 113.470 224.800 ;
        RECT 113.770 224.760 114.470 224.800 ;
        RECT 112.590 224.450 114.470 224.760 ;
        RECT 115.150 224.760 116.230 224.800 ;
        RECT 116.530 224.760 117.400 224.800 ;
        RECT 115.150 224.450 117.400 224.760 ;
        RECT 118.370 224.760 118.990 224.800 ;
        RECT 119.290 224.760 119.950 224.800 ;
        RECT 118.370 224.450 119.950 224.760 ;
        RECT 120.920 224.760 121.750 224.800 ;
        RECT 122.050 224.760 122.710 224.800 ;
        RECT 120.920 224.450 122.710 224.760 ;
        RECT 123.680 224.760 124.510 224.800 ;
        RECT 124.810 224.760 125.400 224.800 ;
        RECT 123.680 224.450 125.400 224.760 ;
        RECT 126.370 224.760 127.270 224.800 ;
        RECT 127.570 224.760 127.705 224.800 ;
        RECT 126.370 224.450 127.705 224.760 ;
        RECT 4.975 220.760 5.325 224.450 ;
        RECT 127.355 224.050 127.705 224.450 ;
        RECT 129.550 224.760 130.030 224.800 ;
        RECT 130.330 224.760 130.660 224.800 ;
        RECT 129.550 224.100 130.660 224.760 ;
        RECT 132.300 224.760 132.790 224.800 ;
        RECT 133.090 224.760 133.550 224.800 ;
        RECT 132.300 224.100 133.550 224.760 ;
        RECT 132.200 223.800 133.550 224.100 ;
        RECT 134.800 224.760 135.550 224.800 ;
        RECT 135.850 224.760 136.350 224.800 ;
        RECT 134.800 223.750 136.350 224.760 ;
        RECT 137.650 224.760 138.310 224.800 ;
        RECT 138.610 224.760 139.150 224.800 ;
        RECT 137.650 223.950 139.150 224.760 ;
        RECT 141.055 224.760 141.070 224.935 ;
        RECT 141.370 224.760 142.160 224.935 ;
        RECT 141.055 224.585 142.160 224.760 ;
        RECT 142.750 224.760 143.830 224.935 ;
        RECT 144.130 224.760 144.600 224.935 ;
        RECT 142.750 224.585 144.600 224.760 ;
        RECT 145.550 224.760 146.590 224.935 ;
        RECT 146.890 224.760 146.935 224.935 ;
        RECT 145.550 224.585 146.935 224.760 ;
        RECT 141.055 223.160 141.405 224.585 ;
        RECT 105.250 144.360 113.830 144.860 ;
        RECT 104.310 142.490 113.830 144.360 ;
        RECT 6.000 141.770 113.830 142.490 ;
        RECT 6.000 138.320 113.250 141.770 ;
        RECT 146.480 140.040 155.490 145.150 ;
        RECT 148.230 139.560 153.090 140.040 ;
        RECT 105.190 136.890 113.250 138.320 ;
        RECT 149.390 9.510 152.030 139.560 ;
        RECT 149.360 5.820 152.950 9.510 ;
        RECT 132.490 1.000 133.390 3.250 ;
        RECT 151.800 1.000 152.720 5.820 ;
        RECT 151.800 0.140 151.810 1.000 ;
        RECT 152.710 0.140 152.720 1.000 ;
  END
END tt_um_r2r_dac
END LIBRARY

