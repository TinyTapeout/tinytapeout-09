module tt_um_urish_giant_ringosc (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \inv_in[0] ;
 wire \inv_in[1000] ;
 wire \inv_in[1001] ;
 wire \inv_in[1002] ;
 wire \inv_in[1003] ;
 wire \inv_in[1004] ;
 wire \inv_in[1005] ;
 wire \inv_in[1006] ;
 wire \inv_in[1007] ;
 wire \inv_in[1008] ;
 wire \inv_in[1009] ;
 wire \inv_in[100] ;
 wire \inv_in[1010] ;
 wire \inv_in[1011] ;
 wire \inv_in[1012] ;
 wire \inv_in[1013] ;
 wire \inv_in[1014] ;
 wire \inv_in[1015] ;
 wire \inv_in[1016] ;
 wire \inv_in[1017] ;
 wire \inv_in[1018] ;
 wire \inv_in[1019] ;
 wire \inv_in[101] ;
 wire \inv_in[1020] ;
 wire \inv_in[1021] ;
 wire \inv_in[1022] ;
 wire \inv_in[1023] ;
 wire \inv_in[1024] ;
 wire \inv_in[1025] ;
 wire \inv_in[1026] ;
 wire \inv_in[1027] ;
 wire \inv_in[1028] ;
 wire \inv_in[1029] ;
 wire \inv_in[102] ;
 wire \inv_in[1030] ;
 wire \inv_in[1031] ;
 wire \inv_in[1032] ;
 wire \inv_in[1033] ;
 wire \inv_in[1034] ;
 wire \inv_in[1035] ;
 wire \inv_in[1036] ;
 wire \inv_in[1037] ;
 wire \inv_in[1038] ;
 wire \inv_in[1039] ;
 wire \inv_in[103] ;
 wire \inv_in[1040] ;
 wire \inv_in[1041] ;
 wire \inv_in[1042] ;
 wire \inv_in[1043] ;
 wire \inv_in[1044] ;
 wire \inv_in[1045] ;
 wire \inv_in[1046] ;
 wire \inv_in[1047] ;
 wire \inv_in[1048] ;
 wire \inv_in[1049] ;
 wire \inv_in[104] ;
 wire \inv_in[1050] ;
 wire \inv_in[1051] ;
 wire \inv_in[1052] ;
 wire \inv_in[1053] ;
 wire \inv_in[1054] ;
 wire \inv_in[1055] ;
 wire \inv_in[1056] ;
 wire \inv_in[1057] ;
 wire \inv_in[1058] ;
 wire \inv_in[1059] ;
 wire \inv_in[105] ;
 wire \inv_in[1060] ;
 wire \inv_in[1061] ;
 wire \inv_in[1062] ;
 wire \inv_in[1063] ;
 wire \inv_in[1064] ;
 wire \inv_in[1065] ;
 wire \inv_in[1066] ;
 wire \inv_in[1067] ;
 wire \inv_in[1068] ;
 wire \inv_in[1069] ;
 wire \inv_in[106] ;
 wire \inv_in[1070] ;
 wire \inv_in[1071] ;
 wire \inv_in[1072] ;
 wire \inv_in[1073] ;
 wire \inv_in[1074] ;
 wire \inv_in[1075] ;
 wire \inv_in[1076] ;
 wire \inv_in[1077] ;
 wire \inv_in[1078] ;
 wire \inv_in[1079] ;
 wire \inv_in[107] ;
 wire \inv_in[1080] ;
 wire \inv_in[1081] ;
 wire \inv_in[1082] ;
 wire \inv_in[1083] ;
 wire \inv_in[1084] ;
 wire \inv_in[1085] ;
 wire \inv_in[1086] ;
 wire \inv_in[1087] ;
 wire \inv_in[1088] ;
 wire \inv_in[1089] ;
 wire \inv_in[108] ;
 wire \inv_in[1090] ;
 wire \inv_in[1091] ;
 wire \inv_in[1092] ;
 wire \inv_in[1093] ;
 wire \inv_in[1094] ;
 wire \inv_in[1095] ;
 wire \inv_in[1096] ;
 wire \inv_in[1097] ;
 wire \inv_in[1098] ;
 wire \inv_in[1099] ;
 wire \inv_in[109] ;
 wire \inv_in[10] ;
 wire \inv_in[1100] ;
 wire \inv_in[1101] ;
 wire \inv_in[1102] ;
 wire \inv_in[1103] ;
 wire \inv_in[1104] ;
 wire \inv_in[1105] ;
 wire \inv_in[1106] ;
 wire \inv_in[1107] ;
 wire \inv_in[1108] ;
 wire \inv_in[1109] ;
 wire \inv_in[110] ;
 wire \inv_in[1110] ;
 wire \inv_in[1111] ;
 wire \inv_in[1112] ;
 wire \inv_in[1113] ;
 wire \inv_in[1114] ;
 wire \inv_in[1115] ;
 wire \inv_in[1116] ;
 wire \inv_in[1117] ;
 wire \inv_in[1118] ;
 wire \inv_in[1119] ;
 wire \inv_in[111] ;
 wire \inv_in[1120] ;
 wire \inv_in[1121] ;
 wire \inv_in[1122] ;
 wire \inv_in[1123] ;
 wire \inv_in[1124] ;
 wire \inv_in[1125] ;
 wire \inv_in[1126] ;
 wire \inv_in[1127] ;
 wire \inv_in[1128] ;
 wire \inv_in[1129] ;
 wire \inv_in[112] ;
 wire \inv_in[1130] ;
 wire \inv_in[1131] ;
 wire \inv_in[1132] ;
 wire \inv_in[1133] ;
 wire \inv_in[1134] ;
 wire \inv_in[1135] ;
 wire \inv_in[1136] ;
 wire \inv_in[1137] ;
 wire \inv_in[1138] ;
 wire \inv_in[1139] ;
 wire \inv_in[113] ;
 wire \inv_in[1140] ;
 wire \inv_in[1141] ;
 wire \inv_in[1142] ;
 wire \inv_in[1143] ;
 wire \inv_in[1144] ;
 wire \inv_in[1145] ;
 wire \inv_in[1146] ;
 wire \inv_in[1147] ;
 wire \inv_in[1148] ;
 wire \inv_in[1149] ;
 wire \inv_in[114] ;
 wire \inv_in[1150] ;
 wire \inv_in[1151] ;
 wire \inv_in[1152] ;
 wire \inv_in[1153] ;
 wire \inv_in[1154] ;
 wire \inv_in[1155] ;
 wire \inv_in[1156] ;
 wire \inv_in[1157] ;
 wire \inv_in[1158] ;
 wire \inv_in[1159] ;
 wire \inv_in[115] ;
 wire \inv_in[1160] ;
 wire \inv_in[1161] ;
 wire \inv_in[1162] ;
 wire \inv_in[1163] ;
 wire \inv_in[1164] ;
 wire \inv_in[1165] ;
 wire \inv_in[1166] ;
 wire \inv_in[1167] ;
 wire \inv_in[1168] ;
 wire \inv_in[1169] ;
 wire \inv_in[116] ;
 wire \inv_in[1170] ;
 wire \inv_in[1171] ;
 wire \inv_in[1172] ;
 wire \inv_in[1173] ;
 wire \inv_in[1174] ;
 wire \inv_in[1175] ;
 wire \inv_in[1176] ;
 wire \inv_in[1177] ;
 wire \inv_in[1178] ;
 wire \inv_in[1179] ;
 wire \inv_in[117] ;
 wire \inv_in[1180] ;
 wire \inv_in[1181] ;
 wire \inv_in[1182] ;
 wire \inv_in[1183] ;
 wire \inv_in[1184] ;
 wire \inv_in[1185] ;
 wire \inv_in[1186] ;
 wire \inv_in[1187] ;
 wire \inv_in[1188] ;
 wire \inv_in[1189] ;
 wire \inv_in[118] ;
 wire \inv_in[1190] ;
 wire \inv_in[1191] ;
 wire \inv_in[1192] ;
 wire \inv_in[1193] ;
 wire \inv_in[1194] ;
 wire \inv_in[1195] ;
 wire \inv_in[1196] ;
 wire \inv_in[1197] ;
 wire \inv_in[1198] ;
 wire \inv_in[1199] ;
 wire \inv_in[119] ;
 wire \inv_in[11] ;
 wire \inv_in[1200] ;
 wire \inv_in[1201] ;
 wire \inv_in[1202] ;
 wire \inv_in[1203] ;
 wire \inv_in[1204] ;
 wire \inv_in[1205] ;
 wire \inv_in[1206] ;
 wire \inv_in[1207] ;
 wire \inv_in[1208] ;
 wire \inv_in[1209] ;
 wire \inv_in[120] ;
 wire \inv_in[1210] ;
 wire \inv_in[1211] ;
 wire \inv_in[1212] ;
 wire \inv_in[1213] ;
 wire \inv_in[1214] ;
 wire \inv_in[1215] ;
 wire \inv_in[1216] ;
 wire \inv_in[1217] ;
 wire \inv_in[1218] ;
 wire \inv_in[1219] ;
 wire \inv_in[121] ;
 wire \inv_in[1220] ;
 wire \inv_in[1221] ;
 wire \inv_in[1222] ;
 wire \inv_in[1223] ;
 wire \inv_in[1224] ;
 wire \inv_in[1225] ;
 wire \inv_in[1226] ;
 wire \inv_in[1227] ;
 wire \inv_in[1228] ;
 wire \inv_in[1229] ;
 wire \inv_in[122] ;
 wire \inv_in[1230] ;
 wire \inv_in[1231] ;
 wire \inv_in[1232] ;
 wire \inv_in[1233] ;
 wire \inv_in[1234] ;
 wire \inv_in[1235] ;
 wire \inv_in[1236] ;
 wire \inv_in[1237] ;
 wire \inv_in[1238] ;
 wire \inv_in[1239] ;
 wire \inv_in[123] ;
 wire \inv_in[1240] ;
 wire \inv_in[1241] ;
 wire \inv_in[1242] ;
 wire \inv_in[1243] ;
 wire \inv_in[1244] ;
 wire \inv_in[1245] ;
 wire \inv_in[1246] ;
 wire \inv_in[1247] ;
 wire \inv_in[1248] ;
 wire \inv_in[1249] ;
 wire \inv_in[124] ;
 wire \inv_in[1250] ;
 wire \inv_in[1251] ;
 wire \inv_in[1252] ;
 wire \inv_in[1253] ;
 wire \inv_in[1254] ;
 wire \inv_in[1255] ;
 wire \inv_in[1256] ;
 wire \inv_in[1257] ;
 wire \inv_in[1258] ;
 wire \inv_in[1259] ;
 wire \inv_in[125] ;
 wire \inv_in[1260] ;
 wire \inv_in[1261] ;
 wire \inv_in[1262] ;
 wire \inv_in[1263] ;
 wire \inv_in[1264] ;
 wire \inv_in[1265] ;
 wire \inv_in[1266] ;
 wire \inv_in[1267] ;
 wire \inv_in[1268] ;
 wire \inv_in[1269] ;
 wire \inv_in[126] ;
 wire \inv_in[1270] ;
 wire \inv_in[1271] ;
 wire \inv_in[1272] ;
 wire \inv_in[1273] ;
 wire \inv_in[1274] ;
 wire \inv_in[1275] ;
 wire \inv_in[1276] ;
 wire \inv_in[1277] ;
 wire \inv_in[1278] ;
 wire \inv_in[1279] ;
 wire \inv_in[127] ;
 wire \inv_in[1280] ;
 wire \inv_in[1281] ;
 wire \inv_in[1282] ;
 wire \inv_in[1283] ;
 wire \inv_in[1284] ;
 wire \inv_in[1285] ;
 wire \inv_in[1286] ;
 wire \inv_in[1287] ;
 wire \inv_in[1288] ;
 wire \inv_in[1289] ;
 wire \inv_in[128] ;
 wire \inv_in[1290] ;
 wire \inv_in[1291] ;
 wire \inv_in[1292] ;
 wire \inv_in[1293] ;
 wire \inv_in[1294] ;
 wire \inv_in[1295] ;
 wire \inv_in[1296] ;
 wire \inv_in[1297] ;
 wire \inv_in[1298] ;
 wire \inv_in[1299] ;
 wire \inv_in[129] ;
 wire \inv_in[12] ;
 wire \inv_in[1300] ;
 wire \inv_in[1301] ;
 wire \inv_in[1302] ;
 wire \inv_in[1303] ;
 wire \inv_in[1304] ;
 wire \inv_in[1305] ;
 wire \inv_in[1306] ;
 wire \inv_in[1307] ;
 wire \inv_in[1308] ;
 wire \inv_in[1309] ;
 wire \inv_in[130] ;
 wire \inv_in[1310] ;
 wire \inv_in[1311] ;
 wire \inv_in[1312] ;
 wire \inv_in[1313] ;
 wire \inv_in[1314] ;
 wire \inv_in[1315] ;
 wire \inv_in[1316] ;
 wire \inv_in[1317] ;
 wire \inv_in[1318] ;
 wire \inv_in[1319] ;
 wire \inv_in[131] ;
 wire \inv_in[1320] ;
 wire \inv_in[1321] ;
 wire \inv_in[1322] ;
 wire \inv_in[1323] ;
 wire \inv_in[1324] ;
 wire \inv_in[1325] ;
 wire \inv_in[1326] ;
 wire \inv_in[1327] ;
 wire \inv_in[1328] ;
 wire \inv_in[1329] ;
 wire \inv_in[132] ;
 wire \inv_in[1330] ;
 wire \inv_in[1331] ;
 wire \inv_in[1332] ;
 wire \inv_in[1333] ;
 wire \inv_in[1334] ;
 wire \inv_in[1335] ;
 wire \inv_in[1336] ;
 wire \inv_in[1337] ;
 wire \inv_in[1338] ;
 wire \inv_in[1339] ;
 wire \inv_in[133] ;
 wire \inv_in[1340] ;
 wire \inv_in[1341] ;
 wire \inv_in[1342] ;
 wire \inv_in[1343] ;
 wire \inv_in[1344] ;
 wire \inv_in[1345] ;
 wire \inv_in[1346] ;
 wire \inv_in[1347] ;
 wire \inv_in[1348] ;
 wire \inv_in[1349] ;
 wire \inv_in[134] ;
 wire \inv_in[1350] ;
 wire \inv_in[1351] ;
 wire \inv_in[1352] ;
 wire \inv_in[1353] ;
 wire \inv_in[1354] ;
 wire \inv_in[1355] ;
 wire \inv_in[1356] ;
 wire \inv_in[1357] ;
 wire \inv_in[1358] ;
 wire \inv_in[1359] ;
 wire \inv_in[135] ;
 wire \inv_in[1360] ;
 wire \inv_in[1361] ;
 wire \inv_in[1362] ;
 wire \inv_in[1363] ;
 wire \inv_in[1364] ;
 wire \inv_in[1365] ;
 wire \inv_in[1366] ;
 wire \inv_in[1367] ;
 wire \inv_in[1368] ;
 wire \inv_in[1369] ;
 wire \inv_in[136] ;
 wire \inv_in[1370] ;
 wire \inv_in[1371] ;
 wire \inv_in[1372] ;
 wire \inv_in[1373] ;
 wire \inv_in[1374] ;
 wire \inv_in[1375] ;
 wire \inv_in[1376] ;
 wire \inv_in[1377] ;
 wire \inv_in[1378] ;
 wire \inv_in[1379] ;
 wire \inv_in[137] ;
 wire \inv_in[1380] ;
 wire \inv_in[1381] ;
 wire \inv_in[1382] ;
 wire \inv_in[1383] ;
 wire \inv_in[1384] ;
 wire \inv_in[1385] ;
 wire \inv_in[1386] ;
 wire \inv_in[1387] ;
 wire \inv_in[1388] ;
 wire \inv_in[1389] ;
 wire \inv_in[138] ;
 wire \inv_in[1390] ;
 wire \inv_in[1391] ;
 wire \inv_in[1392] ;
 wire \inv_in[1393] ;
 wire \inv_in[1394] ;
 wire \inv_in[1395] ;
 wire \inv_in[1396] ;
 wire \inv_in[1397] ;
 wire \inv_in[1398] ;
 wire \inv_in[1399] ;
 wire \inv_in[139] ;
 wire \inv_in[13] ;
 wire \inv_in[1400] ;
 wire \inv_in[1401] ;
 wire \inv_in[1402] ;
 wire \inv_in[1403] ;
 wire \inv_in[1404] ;
 wire \inv_in[1405] ;
 wire \inv_in[1406] ;
 wire \inv_in[1407] ;
 wire \inv_in[1408] ;
 wire \inv_in[1409] ;
 wire \inv_in[140] ;
 wire \inv_in[1410] ;
 wire \inv_in[1411] ;
 wire \inv_in[1412] ;
 wire \inv_in[1413] ;
 wire \inv_in[1414] ;
 wire \inv_in[1415] ;
 wire \inv_in[1416] ;
 wire \inv_in[1417] ;
 wire \inv_in[1418] ;
 wire \inv_in[1419] ;
 wire \inv_in[141] ;
 wire \inv_in[1420] ;
 wire \inv_in[1421] ;
 wire \inv_in[1422] ;
 wire \inv_in[1423] ;
 wire \inv_in[1424] ;
 wire \inv_in[1425] ;
 wire \inv_in[1426] ;
 wire \inv_in[1427] ;
 wire \inv_in[1428] ;
 wire \inv_in[1429] ;
 wire \inv_in[142] ;
 wire \inv_in[1430] ;
 wire \inv_in[1431] ;
 wire \inv_in[1432] ;
 wire \inv_in[1433] ;
 wire \inv_in[1434] ;
 wire \inv_in[1435] ;
 wire \inv_in[1436] ;
 wire \inv_in[1437] ;
 wire \inv_in[1438] ;
 wire \inv_in[1439] ;
 wire \inv_in[143] ;
 wire \inv_in[1440] ;
 wire \inv_in[1441] ;
 wire \inv_in[1442] ;
 wire \inv_in[1443] ;
 wire \inv_in[1444] ;
 wire \inv_in[1445] ;
 wire \inv_in[1446] ;
 wire \inv_in[1447] ;
 wire \inv_in[1448] ;
 wire \inv_in[1449] ;
 wire \inv_in[144] ;
 wire \inv_in[1450] ;
 wire \inv_in[1451] ;
 wire \inv_in[1452] ;
 wire \inv_in[1453] ;
 wire \inv_in[1454] ;
 wire \inv_in[1455] ;
 wire \inv_in[1456] ;
 wire \inv_in[1457] ;
 wire \inv_in[1458] ;
 wire \inv_in[1459] ;
 wire \inv_in[145] ;
 wire \inv_in[1460] ;
 wire \inv_in[1461] ;
 wire \inv_in[1462] ;
 wire \inv_in[1463] ;
 wire \inv_in[1464] ;
 wire \inv_in[1465] ;
 wire \inv_in[1466] ;
 wire \inv_in[1467] ;
 wire \inv_in[1468] ;
 wire \inv_in[1469] ;
 wire \inv_in[146] ;
 wire \inv_in[1470] ;
 wire \inv_in[1471] ;
 wire \inv_in[1472] ;
 wire \inv_in[1473] ;
 wire \inv_in[1474] ;
 wire \inv_in[1475] ;
 wire \inv_in[1476] ;
 wire \inv_in[1477] ;
 wire \inv_in[1478] ;
 wire \inv_in[1479] ;
 wire \inv_in[147] ;
 wire \inv_in[1480] ;
 wire \inv_in[1481] ;
 wire \inv_in[1482] ;
 wire \inv_in[1483] ;
 wire \inv_in[1484] ;
 wire \inv_in[1485] ;
 wire \inv_in[1486] ;
 wire \inv_in[1487] ;
 wire \inv_in[1488] ;
 wire \inv_in[1489] ;
 wire \inv_in[148] ;
 wire \inv_in[1490] ;
 wire \inv_in[1491] ;
 wire \inv_in[1492] ;
 wire \inv_in[1493] ;
 wire \inv_in[1494] ;
 wire \inv_in[1495] ;
 wire \inv_in[1496] ;
 wire \inv_in[1497] ;
 wire \inv_in[1498] ;
 wire \inv_in[1499] ;
 wire \inv_in[149] ;
 wire \inv_in[14] ;
 wire \inv_in[1500] ;
 wire \inv_in[1501] ;
 wire \inv_in[1502] ;
 wire \inv_in[1503] ;
 wire \inv_in[1504] ;
 wire \inv_in[1505] ;
 wire \inv_in[1506] ;
 wire \inv_in[1507] ;
 wire \inv_in[1508] ;
 wire \inv_in[1509] ;
 wire \inv_in[150] ;
 wire \inv_in[1510] ;
 wire \inv_in[1511] ;
 wire \inv_in[1512] ;
 wire \inv_in[1513] ;
 wire \inv_in[1514] ;
 wire \inv_in[1515] ;
 wire \inv_in[1516] ;
 wire \inv_in[1517] ;
 wire \inv_in[1518] ;
 wire \inv_in[1519] ;
 wire \inv_in[151] ;
 wire \inv_in[1520] ;
 wire \inv_in[1521] ;
 wire \inv_in[1522] ;
 wire \inv_in[1523] ;
 wire \inv_in[1524] ;
 wire \inv_in[1525] ;
 wire \inv_in[1526] ;
 wire \inv_in[1527] ;
 wire \inv_in[1528] ;
 wire \inv_in[1529] ;
 wire \inv_in[152] ;
 wire \inv_in[1530] ;
 wire \inv_in[1531] ;
 wire \inv_in[1532] ;
 wire \inv_in[1533] ;
 wire \inv_in[1534] ;
 wire \inv_in[1535] ;
 wire \inv_in[1536] ;
 wire \inv_in[1537] ;
 wire \inv_in[1538] ;
 wire \inv_in[1539] ;
 wire \inv_in[153] ;
 wire \inv_in[1540] ;
 wire \inv_in[1541] ;
 wire \inv_in[1542] ;
 wire \inv_in[1543] ;
 wire \inv_in[1544] ;
 wire \inv_in[1545] ;
 wire \inv_in[1546] ;
 wire \inv_in[1547] ;
 wire \inv_in[1548] ;
 wire \inv_in[1549] ;
 wire \inv_in[154] ;
 wire \inv_in[1550] ;
 wire \inv_in[1551] ;
 wire \inv_in[1552] ;
 wire \inv_in[1553] ;
 wire \inv_in[1554] ;
 wire \inv_in[1555] ;
 wire \inv_in[1556] ;
 wire \inv_in[1557] ;
 wire \inv_in[1558] ;
 wire \inv_in[1559] ;
 wire \inv_in[155] ;
 wire \inv_in[1560] ;
 wire \inv_in[1561] ;
 wire \inv_in[1562] ;
 wire \inv_in[1563] ;
 wire \inv_in[1564] ;
 wire \inv_in[1565] ;
 wire \inv_in[1566] ;
 wire \inv_in[1567] ;
 wire \inv_in[1568] ;
 wire \inv_in[1569] ;
 wire \inv_in[156] ;
 wire \inv_in[1570] ;
 wire \inv_in[1571] ;
 wire \inv_in[1572] ;
 wire \inv_in[1573] ;
 wire \inv_in[1574] ;
 wire \inv_in[1575] ;
 wire \inv_in[1576] ;
 wire \inv_in[1577] ;
 wire \inv_in[1578] ;
 wire \inv_in[1579] ;
 wire \inv_in[157] ;
 wire \inv_in[1580] ;
 wire \inv_in[1581] ;
 wire \inv_in[1582] ;
 wire \inv_in[1583] ;
 wire \inv_in[1584] ;
 wire \inv_in[1585] ;
 wire \inv_in[1586] ;
 wire \inv_in[1587] ;
 wire \inv_in[1588] ;
 wire \inv_in[1589] ;
 wire \inv_in[158] ;
 wire \inv_in[1590] ;
 wire \inv_in[1591] ;
 wire \inv_in[1592] ;
 wire \inv_in[1593] ;
 wire \inv_in[1594] ;
 wire \inv_in[1595] ;
 wire \inv_in[1596] ;
 wire \inv_in[1597] ;
 wire \inv_in[1598] ;
 wire \inv_in[1599] ;
 wire \inv_in[159] ;
 wire \inv_in[15] ;
 wire \inv_in[1600] ;
 wire \inv_in[1601] ;
 wire \inv_in[1602] ;
 wire \inv_in[1603] ;
 wire \inv_in[1604] ;
 wire \inv_in[1605] ;
 wire \inv_in[1606] ;
 wire \inv_in[1607] ;
 wire \inv_in[1608] ;
 wire \inv_in[1609] ;
 wire \inv_in[160] ;
 wire \inv_in[1610] ;
 wire \inv_in[1611] ;
 wire \inv_in[1612] ;
 wire \inv_in[1613] ;
 wire \inv_in[1614] ;
 wire \inv_in[1615] ;
 wire \inv_in[1616] ;
 wire \inv_in[1617] ;
 wire \inv_in[1618] ;
 wire \inv_in[1619] ;
 wire \inv_in[161] ;
 wire \inv_in[1620] ;
 wire \inv_in[1621] ;
 wire \inv_in[1622] ;
 wire \inv_in[1623] ;
 wire \inv_in[1624] ;
 wire \inv_in[1625] ;
 wire \inv_in[1626] ;
 wire \inv_in[1627] ;
 wire \inv_in[1628] ;
 wire \inv_in[1629] ;
 wire \inv_in[162] ;
 wire \inv_in[1630] ;
 wire \inv_in[1631] ;
 wire \inv_in[1632] ;
 wire \inv_in[1633] ;
 wire \inv_in[1634] ;
 wire \inv_in[1635] ;
 wire \inv_in[1636] ;
 wire \inv_in[1637] ;
 wire \inv_in[1638] ;
 wire \inv_in[1639] ;
 wire \inv_in[163] ;
 wire \inv_in[1640] ;
 wire \inv_in[1641] ;
 wire \inv_in[1642] ;
 wire \inv_in[1643] ;
 wire \inv_in[1644] ;
 wire \inv_in[1645] ;
 wire \inv_in[1646] ;
 wire \inv_in[1647] ;
 wire \inv_in[1648] ;
 wire \inv_in[1649] ;
 wire \inv_in[164] ;
 wire \inv_in[1650] ;
 wire \inv_in[1651] ;
 wire \inv_in[1652] ;
 wire \inv_in[1653] ;
 wire \inv_in[1654] ;
 wire \inv_in[1655] ;
 wire \inv_in[1656] ;
 wire \inv_in[1657] ;
 wire \inv_in[1658] ;
 wire \inv_in[1659] ;
 wire \inv_in[165] ;
 wire \inv_in[1660] ;
 wire \inv_in[1661] ;
 wire \inv_in[1662] ;
 wire \inv_in[1663] ;
 wire \inv_in[1664] ;
 wire \inv_in[1665] ;
 wire \inv_in[1666] ;
 wire \inv_in[1667] ;
 wire \inv_in[1668] ;
 wire \inv_in[1669] ;
 wire \inv_in[166] ;
 wire \inv_in[1670] ;
 wire \inv_in[1671] ;
 wire \inv_in[1672] ;
 wire \inv_in[1673] ;
 wire \inv_in[1674] ;
 wire \inv_in[1675] ;
 wire \inv_in[1676] ;
 wire \inv_in[1677] ;
 wire \inv_in[1678] ;
 wire \inv_in[1679] ;
 wire \inv_in[167] ;
 wire \inv_in[1680] ;
 wire \inv_in[1681] ;
 wire \inv_in[1682] ;
 wire \inv_in[1683] ;
 wire \inv_in[1684] ;
 wire \inv_in[1685] ;
 wire \inv_in[1686] ;
 wire \inv_in[1687] ;
 wire \inv_in[1688] ;
 wire \inv_in[1689] ;
 wire \inv_in[168] ;
 wire \inv_in[1690] ;
 wire \inv_in[1691] ;
 wire \inv_in[1692] ;
 wire \inv_in[1693] ;
 wire \inv_in[1694] ;
 wire \inv_in[1695] ;
 wire \inv_in[1696] ;
 wire \inv_in[1697] ;
 wire \inv_in[1698] ;
 wire \inv_in[1699] ;
 wire \inv_in[169] ;
 wire \inv_in[16] ;
 wire \inv_in[1700] ;
 wire \inv_in[1701] ;
 wire \inv_in[1702] ;
 wire \inv_in[1703] ;
 wire \inv_in[1704] ;
 wire \inv_in[1705] ;
 wire \inv_in[1706] ;
 wire \inv_in[1707] ;
 wire \inv_in[1708] ;
 wire \inv_in[1709] ;
 wire \inv_in[170] ;
 wire \inv_in[1710] ;
 wire \inv_in[1711] ;
 wire \inv_in[1712] ;
 wire \inv_in[1713] ;
 wire \inv_in[1714] ;
 wire \inv_in[1715] ;
 wire \inv_in[1716] ;
 wire \inv_in[1717] ;
 wire \inv_in[1718] ;
 wire \inv_in[1719] ;
 wire \inv_in[171] ;
 wire \inv_in[1720] ;
 wire \inv_in[1721] ;
 wire \inv_in[1722] ;
 wire \inv_in[1723] ;
 wire \inv_in[1724] ;
 wire \inv_in[1725] ;
 wire \inv_in[1726] ;
 wire \inv_in[1727] ;
 wire \inv_in[1728] ;
 wire \inv_in[1729] ;
 wire \inv_in[172] ;
 wire \inv_in[1730] ;
 wire \inv_in[1731] ;
 wire \inv_in[1732] ;
 wire \inv_in[1733] ;
 wire \inv_in[1734] ;
 wire \inv_in[1735] ;
 wire \inv_in[1736] ;
 wire \inv_in[1737] ;
 wire \inv_in[1738] ;
 wire \inv_in[1739] ;
 wire \inv_in[173] ;
 wire \inv_in[1740] ;
 wire \inv_in[1741] ;
 wire \inv_in[1742] ;
 wire \inv_in[1743] ;
 wire \inv_in[1744] ;
 wire \inv_in[1745] ;
 wire \inv_in[1746] ;
 wire \inv_in[1747] ;
 wire \inv_in[1748] ;
 wire \inv_in[1749] ;
 wire \inv_in[174] ;
 wire \inv_in[1750] ;
 wire \inv_in[1751] ;
 wire \inv_in[1752] ;
 wire \inv_in[1753] ;
 wire \inv_in[1754] ;
 wire \inv_in[1755] ;
 wire \inv_in[1756] ;
 wire \inv_in[1757] ;
 wire \inv_in[1758] ;
 wire \inv_in[1759] ;
 wire \inv_in[175] ;
 wire \inv_in[1760] ;
 wire \inv_in[1761] ;
 wire \inv_in[1762] ;
 wire \inv_in[1763] ;
 wire \inv_in[1764] ;
 wire \inv_in[1765] ;
 wire \inv_in[1766] ;
 wire \inv_in[1767] ;
 wire \inv_in[1768] ;
 wire \inv_in[1769] ;
 wire \inv_in[176] ;
 wire \inv_in[1770] ;
 wire \inv_in[1771] ;
 wire \inv_in[1772] ;
 wire \inv_in[1773] ;
 wire \inv_in[1774] ;
 wire \inv_in[1775] ;
 wire \inv_in[1776] ;
 wire \inv_in[1777] ;
 wire \inv_in[1778] ;
 wire \inv_in[1779] ;
 wire \inv_in[177] ;
 wire \inv_in[1780] ;
 wire \inv_in[1781] ;
 wire \inv_in[1782] ;
 wire \inv_in[1783] ;
 wire \inv_in[1784] ;
 wire \inv_in[1785] ;
 wire \inv_in[1786] ;
 wire \inv_in[1787] ;
 wire \inv_in[1788] ;
 wire \inv_in[1789] ;
 wire \inv_in[178] ;
 wire \inv_in[1790] ;
 wire \inv_in[1791] ;
 wire \inv_in[1792] ;
 wire \inv_in[1793] ;
 wire \inv_in[1794] ;
 wire \inv_in[1795] ;
 wire \inv_in[1796] ;
 wire \inv_in[1797] ;
 wire \inv_in[1798] ;
 wire \inv_in[1799] ;
 wire \inv_in[179] ;
 wire \inv_in[17] ;
 wire \inv_in[1800] ;
 wire \inv_in[1801] ;
 wire \inv_in[1802] ;
 wire \inv_in[1803] ;
 wire \inv_in[1804] ;
 wire \inv_in[1805] ;
 wire \inv_in[1806] ;
 wire \inv_in[1807] ;
 wire \inv_in[1808] ;
 wire \inv_in[1809] ;
 wire \inv_in[180] ;
 wire \inv_in[1810] ;
 wire \inv_in[1811] ;
 wire \inv_in[1812] ;
 wire \inv_in[1813] ;
 wire \inv_in[1814] ;
 wire \inv_in[1815] ;
 wire \inv_in[1816] ;
 wire \inv_in[1817] ;
 wire \inv_in[1818] ;
 wire \inv_in[1819] ;
 wire \inv_in[181] ;
 wire \inv_in[1820] ;
 wire \inv_in[1821] ;
 wire \inv_in[1822] ;
 wire \inv_in[1823] ;
 wire \inv_in[1824] ;
 wire \inv_in[1825] ;
 wire \inv_in[1826] ;
 wire \inv_in[1827] ;
 wire \inv_in[1828] ;
 wire \inv_in[1829] ;
 wire \inv_in[182] ;
 wire \inv_in[1830] ;
 wire \inv_in[1831] ;
 wire \inv_in[1832] ;
 wire \inv_in[1833] ;
 wire \inv_in[1834] ;
 wire \inv_in[1835] ;
 wire \inv_in[1836] ;
 wire \inv_in[1837] ;
 wire \inv_in[1838] ;
 wire \inv_in[1839] ;
 wire \inv_in[183] ;
 wire \inv_in[1840] ;
 wire \inv_in[1841] ;
 wire \inv_in[1842] ;
 wire \inv_in[1843] ;
 wire \inv_in[1844] ;
 wire \inv_in[1845] ;
 wire \inv_in[1846] ;
 wire \inv_in[1847] ;
 wire \inv_in[1848] ;
 wire \inv_in[1849] ;
 wire \inv_in[184] ;
 wire \inv_in[1850] ;
 wire \inv_in[1851] ;
 wire \inv_in[1852] ;
 wire \inv_in[1853] ;
 wire \inv_in[1854] ;
 wire \inv_in[1855] ;
 wire \inv_in[1856] ;
 wire \inv_in[1857] ;
 wire \inv_in[1858] ;
 wire \inv_in[1859] ;
 wire \inv_in[185] ;
 wire \inv_in[1860] ;
 wire \inv_in[1861] ;
 wire \inv_in[1862] ;
 wire \inv_in[1863] ;
 wire \inv_in[1864] ;
 wire \inv_in[1865] ;
 wire \inv_in[1866] ;
 wire \inv_in[1867] ;
 wire \inv_in[1868] ;
 wire \inv_in[1869] ;
 wire \inv_in[186] ;
 wire \inv_in[1870] ;
 wire \inv_in[1871] ;
 wire \inv_in[1872] ;
 wire \inv_in[1873] ;
 wire \inv_in[1874] ;
 wire \inv_in[1875] ;
 wire \inv_in[1876] ;
 wire \inv_in[1877] ;
 wire \inv_in[1878] ;
 wire \inv_in[1879] ;
 wire \inv_in[187] ;
 wire \inv_in[1880] ;
 wire \inv_in[1881] ;
 wire \inv_in[1882] ;
 wire \inv_in[1883] ;
 wire \inv_in[1884] ;
 wire \inv_in[1885] ;
 wire \inv_in[1886] ;
 wire \inv_in[1887] ;
 wire \inv_in[1888] ;
 wire \inv_in[1889] ;
 wire \inv_in[188] ;
 wire \inv_in[1890] ;
 wire \inv_in[1891] ;
 wire \inv_in[1892] ;
 wire \inv_in[1893] ;
 wire \inv_in[1894] ;
 wire \inv_in[1895] ;
 wire \inv_in[1896] ;
 wire \inv_in[1897] ;
 wire \inv_in[1898] ;
 wire \inv_in[1899] ;
 wire \inv_in[189] ;
 wire \inv_in[18] ;
 wire \inv_in[1900] ;
 wire \inv_in[1901] ;
 wire \inv_in[1902] ;
 wire \inv_in[1903] ;
 wire \inv_in[1904] ;
 wire \inv_in[1905] ;
 wire \inv_in[1906] ;
 wire \inv_in[1907] ;
 wire \inv_in[1908] ;
 wire \inv_in[1909] ;
 wire \inv_in[190] ;
 wire \inv_in[1910] ;
 wire \inv_in[1911] ;
 wire \inv_in[1912] ;
 wire \inv_in[1913] ;
 wire \inv_in[1914] ;
 wire \inv_in[1915] ;
 wire \inv_in[1916] ;
 wire \inv_in[1917] ;
 wire \inv_in[1918] ;
 wire \inv_in[1919] ;
 wire \inv_in[191] ;
 wire \inv_in[1920] ;
 wire \inv_in[1921] ;
 wire \inv_in[1922] ;
 wire \inv_in[1923] ;
 wire \inv_in[1924] ;
 wire \inv_in[1925] ;
 wire \inv_in[1926] ;
 wire \inv_in[1927] ;
 wire \inv_in[1928] ;
 wire \inv_in[1929] ;
 wire \inv_in[192] ;
 wire \inv_in[1930] ;
 wire \inv_in[1931] ;
 wire \inv_in[1932] ;
 wire \inv_in[1933] ;
 wire \inv_in[1934] ;
 wire \inv_in[1935] ;
 wire \inv_in[1936] ;
 wire \inv_in[1937] ;
 wire \inv_in[1938] ;
 wire \inv_in[1939] ;
 wire \inv_in[193] ;
 wire \inv_in[1940] ;
 wire \inv_in[1941] ;
 wire \inv_in[1942] ;
 wire \inv_in[1943] ;
 wire \inv_in[1944] ;
 wire \inv_in[1945] ;
 wire \inv_in[1946] ;
 wire \inv_in[1947] ;
 wire \inv_in[1948] ;
 wire \inv_in[1949] ;
 wire \inv_in[194] ;
 wire \inv_in[1950] ;
 wire \inv_in[1951] ;
 wire \inv_in[1952] ;
 wire \inv_in[1953] ;
 wire \inv_in[1954] ;
 wire \inv_in[1955] ;
 wire \inv_in[1956] ;
 wire \inv_in[1957] ;
 wire \inv_in[1958] ;
 wire \inv_in[1959] ;
 wire \inv_in[195] ;
 wire \inv_in[1960] ;
 wire \inv_in[1961] ;
 wire \inv_in[1962] ;
 wire \inv_in[1963] ;
 wire \inv_in[1964] ;
 wire \inv_in[1965] ;
 wire \inv_in[1966] ;
 wire \inv_in[1967] ;
 wire \inv_in[1968] ;
 wire \inv_in[1969] ;
 wire \inv_in[196] ;
 wire \inv_in[1970] ;
 wire \inv_in[1971] ;
 wire \inv_in[1972] ;
 wire \inv_in[1973] ;
 wire \inv_in[1974] ;
 wire \inv_in[1975] ;
 wire \inv_in[1976] ;
 wire \inv_in[1977] ;
 wire \inv_in[1978] ;
 wire \inv_in[1979] ;
 wire \inv_in[197] ;
 wire \inv_in[1980] ;
 wire \inv_in[1981] ;
 wire \inv_in[1982] ;
 wire \inv_in[1983] ;
 wire \inv_in[1984] ;
 wire \inv_in[1985] ;
 wire \inv_in[1986] ;
 wire \inv_in[1987] ;
 wire \inv_in[1988] ;
 wire \inv_in[1989] ;
 wire \inv_in[198] ;
 wire \inv_in[1990] ;
 wire \inv_in[1991] ;
 wire \inv_in[1992] ;
 wire \inv_in[1993] ;
 wire \inv_in[1994] ;
 wire \inv_in[1995] ;
 wire \inv_in[1996] ;
 wire \inv_in[1997] ;
 wire \inv_in[1998] ;
 wire \inv_in[1999] ;
 wire \inv_in[199] ;
 wire \inv_in[19] ;
 wire \inv_in[1] ;
 wire \inv_in[2000] ;
 wire \inv_in[2001] ;
 wire \inv_in[2002] ;
 wire \inv_in[2003] ;
 wire \inv_in[2004] ;
 wire \inv_in[2005] ;
 wire \inv_in[2006] ;
 wire \inv_in[2007] ;
 wire \inv_in[2008] ;
 wire \inv_in[2009] ;
 wire \inv_in[200] ;
 wire \inv_in[2010] ;
 wire \inv_in[2011] ;
 wire \inv_in[2012] ;
 wire \inv_in[2013] ;
 wire \inv_in[2014] ;
 wire \inv_in[2015] ;
 wire \inv_in[2016] ;
 wire \inv_in[2017] ;
 wire \inv_in[2018] ;
 wire \inv_in[2019] ;
 wire \inv_in[201] ;
 wire \inv_in[2020] ;
 wire \inv_in[2021] ;
 wire \inv_in[2022] ;
 wire \inv_in[2023] ;
 wire \inv_in[2024] ;
 wire \inv_in[2025] ;
 wire \inv_in[2026] ;
 wire \inv_in[2027] ;
 wire \inv_in[2028] ;
 wire \inv_in[2029] ;
 wire \inv_in[202] ;
 wire \inv_in[2030] ;
 wire \inv_in[2031] ;
 wire \inv_in[2032] ;
 wire \inv_in[2033] ;
 wire \inv_in[2034] ;
 wire \inv_in[2035] ;
 wire \inv_in[2036] ;
 wire \inv_in[2037] ;
 wire \inv_in[2038] ;
 wire \inv_in[2039] ;
 wire \inv_in[203] ;
 wire \inv_in[2040] ;
 wire \inv_in[2041] ;
 wire \inv_in[2042] ;
 wire \inv_in[2043] ;
 wire \inv_in[2044] ;
 wire \inv_in[2045] ;
 wire \inv_in[2046] ;
 wire \inv_in[2047] ;
 wire \inv_in[2048] ;
 wire \inv_in[2049] ;
 wire \inv_in[204] ;
 wire \inv_in[2050] ;
 wire \inv_in[2051] ;
 wire \inv_in[2052] ;
 wire \inv_in[2053] ;
 wire \inv_in[2054] ;
 wire \inv_in[2055] ;
 wire \inv_in[2056] ;
 wire \inv_in[2057] ;
 wire \inv_in[2058] ;
 wire \inv_in[2059] ;
 wire \inv_in[205] ;
 wire \inv_in[2060] ;
 wire \inv_in[2061] ;
 wire \inv_in[2062] ;
 wire \inv_in[2063] ;
 wire \inv_in[2064] ;
 wire \inv_in[2065] ;
 wire \inv_in[2066] ;
 wire \inv_in[2067] ;
 wire \inv_in[2068] ;
 wire \inv_in[2069] ;
 wire \inv_in[206] ;
 wire \inv_in[2070] ;
 wire \inv_in[2071] ;
 wire \inv_in[2072] ;
 wire \inv_in[2073] ;
 wire \inv_in[2074] ;
 wire \inv_in[2075] ;
 wire \inv_in[2076] ;
 wire \inv_in[2077] ;
 wire \inv_in[2078] ;
 wire \inv_in[2079] ;
 wire \inv_in[207] ;
 wire \inv_in[2080] ;
 wire \inv_in[2081] ;
 wire \inv_in[2082] ;
 wire \inv_in[2083] ;
 wire \inv_in[2084] ;
 wire \inv_in[2085] ;
 wire \inv_in[2086] ;
 wire \inv_in[2087] ;
 wire \inv_in[2088] ;
 wire \inv_in[2089] ;
 wire \inv_in[208] ;
 wire \inv_in[2090] ;
 wire \inv_in[2091] ;
 wire \inv_in[2092] ;
 wire \inv_in[2093] ;
 wire \inv_in[2094] ;
 wire \inv_in[2095] ;
 wire \inv_in[2096] ;
 wire \inv_in[2097] ;
 wire \inv_in[2098] ;
 wire \inv_in[2099] ;
 wire \inv_in[209] ;
 wire \inv_in[20] ;
 wire \inv_in[2100] ;
 wire \inv_in[2101] ;
 wire \inv_in[2102] ;
 wire \inv_in[2103] ;
 wire \inv_in[2104] ;
 wire \inv_in[2105] ;
 wire \inv_in[2106] ;
 wire \inv_in[2107] ;
 wire \inv_in[2108] ;
 wire \inv_in[2109] ;
 wire \inv_in[210] ;
 wire \inv_in[2110] ;
 wire \inv_in[2111] ;
 wire \inv_in[2112] ;
 wire \inv_in[2113] ;
 wire \inv_in[2114] ;
 wire \inv_in[2115] ;
 wire \inv_in[2116] ;
 wire \inv_in[2117] ;
 wire \inv_in[2118] ;
 wire \inv_in[2119] ;
 wire \inv_in[211] ;
 wire \inv_in[2120] ;
 wire \inv_in[2121] ;
 wire \inv_in[2122] ;
 wire \inv_in[2123] ;
 wire \inv_in[2124] ;
 wire \inv_in[2125] ;
 wire \inv_in[2126] ;
 wire \inv_in[2127] ;
 wire \inv_in[2128] ;
 wire \inv_in[2129] ;
 wire \inv_in[212] ;
 wire \inv_in[2130] ;
 wire \inv_in[2131] ;
 wire \inv_in[2132] ;
 wire \inv_in[2133] ;
 wire \inv_in[2134] ;
 wire \inv_in[2135] ;
 wire \inv_in[2136] ;
 wire \inv_in[2137] ;
 wire \inv_in[2138] ;
 wire \inv_in[2139] ;
 wire \inv_in[213] ;
 wire \inv_in[2140] ;
 wire \inv_in[2141] ;
 wire \inv_in[2142] ;
 wire \inv_in[2143] ;
 wire \inv_in[2144] ;
 wire \inv_in[2145] ;
 wire \inv_in[2146] ;
 wire \inv_in[2147] ;
 wire \inv_in[2148] ;
 wire \inv_in[2149] ;
 wire \inv_in[214] ;
 wire \inv_in[2150] ;
 wire \inv_in[2151] ;
 wire \inv_in[2152] ;
 wire \inv_in[2153] ;
 wire \inv_in[2154] ;
 wire \inv_in[2155] ;
 wire \inv_in[2156] ;
 wire \inv_in[2157] ;
 wire \inv_in[2158] ;
 wire \inv_in[2159] ;
 wire \inv_in[215] ;
 wire \inv_in[2160] ;
 wire \inv_in[2161] ;
 wire \inv_in[2162] ;
 wire \inv_in[2163] ;
 wire \inv_in[2164] ;
 wire \inv_in[2165] ;
 wire \inv_in[2166] ;
 wire \inv_in[2167] ;
 wire \inv_in[2168] ;
 wire \inv_in[2169] ;
 wire \inv_in[216] ;
 wire \inv_in[2170] ;
 wire \inv_in[2171] ;
 wire \inv_in[2172] ;
 wire \inv_in[2173] ;
 wire \inv_in[2174] ;
 wire \inv_in[2175] ;
 wire \inv_in[2176] ;
 wire \inv_in[2177] ;
 wire \inv_in[2178] ;
 wire \inv_in[2179] ;
 wire \inv_in[217] ;
 wire \inv_in[2180] ;
 wire \inv_in[2181] ;
 wire \inv_in[2182] ;
 wire \inv_in[2183] ;
 wire \inv_in[2184] ;
 wire \inv_in[2185] ;
 wire \inv_in[2186] ;
 wire \inv_in[2187] ;
 wire \inv_in[2188] ;
 wire \inv_in[2189] ;
 wire \inv_in[218] ;
 wire \inv_in[2190] ;
 wire \inv_in[2191] ;
 wire \inv_in[2192] ;
 wire \inv_in[2193] ;
 wire \inv_in[2194] ;
 wire \inv_in[2195] ;
 wire \inv_in[2196] ;
 wire \inv_in[2197] ;
 wire \inv_in[2198] ;
 wire \inv_in[2199] ;
 wire \inv_in[219] ;
 wire \inv_in[21] ;
 wire \inv_in[2200] ;
 wire \inv_in[2201] ;
 wire \inv_in[2202] ;
 wire \inv_in[2203] ;
 wire \inv_in[2204] ;
 wire \inv_in[2205] ;
 wire \inv_in[2206] ;
 wire \inv_in[2207] ;
 wire \inv_in[2208] ;
 wire \inv_in[2209] ;
 wire \inv_in[220] ;
 wire \inv_in[2210] ;
 wire \inv_in[2211] ;
 wire \inv_in[2212] ;
 wire \inv_in[2213] ;
 wire \inv_in[2214] ;
 wire \inv_in[2215] ;
 wire \inv_in[2216] ;
 wire \inv_in[2217] ;
 wire \inv_in[2218] ;
 wire \inv_in[2219] ;
 wire \inv_in[221] ;
 wire \inv_in[2220] ;
 wire \inv_in[2221] ;
 wire \inv_in[2222] ;
 wire \inv_in[2223] ;
 wire \inv_in[2224] ;
 wire \inv_in[2225] ;
 wire \inv_in[2226] ;
 wire \inv_in[2227] ;
 wire \inv_in[2228] ;
 wire \inv_in[2229] ;
 wire \inv_in[222] ;
 wire \inv_in[2230] ;
 wire \inv_in[2231] ;
 wire \inv_in[2232] ;
 wire \inv_in[2233] ;
 wire \inv_in[2234] ;
 wire \inv_in[2235] ;
 wire \inv_in[2236] ;
 wire \inv_in[2237] ;
 wire \inv_in[2238] ;
 wire \inv_in[2239] ;
 wire \inv_in[223] ;
 wire \inv_in[2240] ;
 wire \inv_in[2241] ;
 wire \inv_in[2242] ;
 wire \inv_in[2243] ;
 wire \inv_in[2244] ;
 wire \inv_in[2245] ;
 wire \inv_in[2246] ;
 wire \inv_in[2247] ;
 wire \inv_in[2248] ;
 wire \inv_in[2249] ;
 wire \inv_in[224] ;
 wire \inv_in[2250] ;
 wire \inv_in[2251] ;
 wire \inv_in[2252] ;
 wire \inv_in[2253] ;
 wire \inv_in[2254] ;
 wire \inv_in[2255] ;
 wire \inv_in[2256] ;
 wire \inv_in[2257] ;
 wire \inv_in[2258] ;
 wire \inv_in[2259] ;
 wire \inv_in[225] ;
 wire \inv_in[2260] ;
 wire \inv_in[2261] ;
 wire \inv_in[2262] ;
 wire \inv_in[2263] ;
 wire \inv_in[2264] ;
 wire \inv_in[2265] ;
 wire \inv_in[2266] ;
 wire \inv_in[2267] ;
 wire \inv_in[2268] ;
 wire \inv_in[2269] ;
 wire \inv_in[226] ;
 wire \inv_in[2270] ;
 wire \inv_in[2271] ;
 wire \inv_in[2272] ;
 wire \inv_in[2273] ;
 wire \inv_in[2274] ;
 wire \inv_in[2275] ;
 wire \inv_in[2276] ;
 wire \inv_in[2277] ;
 wire \inv_in[2278] ;
 wire \inv_in[2279] ;
 wire \inv_in[227] ;
 wire \inv_in[2280] ;
 wire \inv_in[2281] ;
 wire \inv_in[2282] ;
 wire \inv_in[2283] ;
 wire \inv_in[2284] ;
 wire \inv_in[2285] ;
 wire \inv_in[2286] ;
 wire \inv_in[2287] ;
 wire \inv_in[2288] ;
 wire \inv_in[2289] ;
 wire \inv_in[228] ;
 wire \inv_in[2290] ;
 wire \inv_in[2291] ;
 wire \inv_in[2292] ;
 wire \inv_in[2293] ;
 wire \inv_in[2294] ;
 wire \inv_in[2295] ;
 wire \inv_in[2296] ;
 wire \inv_in[2297] ;
 wire \inv_in[2298] ;
 wire \inv_in[2299] ;
 wire \inv_in[229] ;
 wire \inv_in[22] ;
 wire \inv_in[2300] ;
 wire \inv_in[2301] ;
 wire \inv_in[2302] ;
 wire \inv_in[2303] ;
 wire \inv_in[2304] ;
 wire \inv_in[2305] ;
 wire \inv_in[2306] ;
 wire \inv_in[2307] ;
 wire \inv_in[2308] ;
 wire \inv_in[2309] ;
 wire \inv_in[230] ;
 wire \inv_in[2310] ;
 wire \inv_in[2311] ;
 wire \inv_in[2312] ;
 wire \inv_in[2313] ;
 wire \inv_in[2314] ;
 wire \inv_in[2315] ;
 wire \inv_in[2316] ;
 wire \inv_in[2317] ;
 wire \inv_in[2318] ;
 wire \inv_in[2319] ;
 wire \inv_in[231] ;
 wire \inv_in[2320] ;
 wire \inv_in[2321] ;
 wire \inv_in[2322] ;
 wire \inv_in[2323] ;
 wire \inv_in[2324] ;
 wire \inv_in[2325] ;
 wire \inv_in[2326] ;
 wire \inv_in[2327] ;
 wire \inv_in[2328] ;
 wire \inv_in[2329] ;
 wire \inv_in[232] ;
 wire \inv_in[2330] ;
 wire \inv_in[2331] ;
 wire \inv_in[2332] ;
 wire \inv_in[2333] ;
 wire \inv_in[2334] ;
 wire \inv_in[2335] ;
 wire \inv_in[2336] ;
 wire \inv_in[2337] ;
 wire \inv_in[2338] ;
 wire \inv_in[2339] ;
 wire \inv_in[233] ;
 wire \inv_in[2340] ;
 wire \inv_in[2341] ;
 wire \inv_in[2342] ;
 wire \inv_in[2343] ;
 wire \inv_in[2344] ;
 wire \inv_in[2345] ;
 wire \inv_in[2346] ;
 wire \inv_in[2347] ;
 wire \inv_in[2348] ;
 wire \inv_in[2349] ;
 wire \inv_in[234] ;
 wire \inv_in[2350] ;
 wire \inv_in[2351] ;
 wire \inv_in[2352] ;
 wire \inv_in[2353] ;
 wire \inv_in[2354] ;
 wire \inv_in[2355] ;
 wire \inv_in[2356] ;
 wire \inv_in[2357] ;
 wire \inv_in[2358] ;
 wire \inv_in[2359] ;
 wire \inv_in[235] ;
 wire \inv_in[2360] ;
 wire \inv_in[2361] ;
 wire \inv_in[2362] ;
 wire \inv_in[2363] ;
 wire \inv_in[2364] ;
 wire \inv_in[2365] ;
 wire \inv_in[2366] ;
 wire \inv_in[2367] ;
 wire \inv_in[2368] ;
 wire \inv_in[2369] ;
 wire \inv_in[236] ;
 wire \inv_in[2370] ;
 wire \inv_in[2371] ;
 wire \inv_in[2372] ;
 wire \inv_in[2373] ;
 wire \inv_in[2374] ;
 wire \inv_in[2375] ;
 wire \inv_in[2376] ;
 wire \inv_in[2377] ;
 wire \inv_in[2378] ;
 wire \inv_in[2379] ;
 wire \inv_in[237] ;
 wire \inv_in[2380] ;
 wire \inv_in[2381] ;
 wire \inv_in[2382] ;
 wire \inv_in[2383] ;
 wire \inv_in[2384] ;
 wire \inv_in[2385] ;
 wire \inv_in[2386] ;
 wire \inv_in[2387] ;
 wire \inv_in[2388] ;
 wire \inv_in[2389] ;
 wire \inv_in[238] ;
 wire \inv_in[2390] ;
 wire \inv_in[2391] ;
 wire \inv_in[2392] ;
 wire \inv_in[2393] ;
 wire \inv_in[2394] ;
 wire \inv_in[2395] ;
 wire \inv_in[2396] ;
 wire \inv_in[2397] ;
 wire \inv_in[2398] ;
 wire \inv_in[2399] ;
 wire \inv_in[239] ;
 wire \inv_in[23] ;
 wire \inv_in[2400] ;
 wire \inv_in[2401] ;
 wire \inv_in[2402] ;
 wire \inv_in[2403] ;
 wire \inv_in[2404] ;
 wire \inv_in[2405] ;
 wire \inv_in[2406] ;
 wire \inv_in[2407] ;
 wire \inv_in[2408] ;
 wire \inv_in[2409] ;
 wire \inv_in[240] ;
 wire \inv_in[2410] ;
 wire \inv_in[2411] ;
 wire \inv_in[2412] ;
 wire \inv_in[2413] ;
 wire \inv_in[2414] ;
 wire \inv_in[2415] ;
 wire \inv_in[2416] ;
 wire \inv_in[2417] ;
 wire \inv_in[2418] ;
 wire \inv_in[2419] ;
 wire \inv_in[241] ;
 wire \inv_in[2420] ;
 wire \inv_in[2421] ;
 wire \inv_in[2422] ;
 wire \inv_in[2423] ;
 wire \inv_in[2424] ;
 wire \inv_in[2425] ;
 wire \inv_in[2426] ;
 wire \inv_in[2427] ;
 wire \inv_in[2428] ;
 wire \inv_in[2429] ;
 wire \inv_in[242] ;
 wire \inv_in[2430] ;
 wire \inv_in[2431] ;
 wire \inv_in[2432] ;
 wire \inv_in[2433] ;
 wire \inv_in[2434] ;
 wire \inv_in[2435] ;
 wire \inv_in[2436] ;
 wire \inv_in[2437] ;
 wire \inv_in[2438] ;
 wire \inv_in[2439] ;
 wire \inv_in[243] ;
 wire \inv_in[2440] ;
 wire \inv_in[2441] ;
 wire \inv_in[2442] ;
 wire \inv_in[2443] ;
 wire \inv_in[2444] ;
 wire \inv_in[2445] ;
 wire \inv_in[2446] ;
 wire \inv_in[2447] ;
 wire \inv_in[2448] ;
 wire \inv_in[2449] ;
 wire \inv_in[244] ;
 wire \inv_in[2450] ;
 wire \inv_in[2451] ;
 wire \inv_in[2452] ;
 wire \inv_in[2453] ;
 wire \inv_in[2454] ;
 wire \inv_in[2455] ;
 wire \inv_in[2456] ;
 wire \inv_in[2457] ;
 wire \inv_in[2458] ;
 wire \inv_in[2459] ;
 wire \inv_in[245] ;
 wire \inv_in[2460] ;
 wire \inv_in[2461] ;
 wire \inv_in[2462] ;
 wire \inv_in[2463] ;
 wire \inv_in[2464] ;
 wire \inv_in[2465] ;
 wire \inv_in[2466] ;
 wire \inv_in[2467] ;
 wire \inv_in[2468] ;
 wire \inv_in[2469] ;
 wire \inv_in[246] ;
 wire \inv_in[2470] ;
 wire \inv_in[2471] ;
 wire \inv_in[2472] ;
 wire \inv_in[2473] ;
 wire \inv_in[2474] ;
 wire \inv_in[2475] ;
 wire \inv_in[2476] ;
 wire \inv_in[2477] ;
 wire \inv_in[2478] ;
 wire \inv_in[2479] ;
 wire \inv_in[247] ;
 wire \inv_in[2480] ;
 wire \inv_in[2481] ;
 wire \inv_in[2482] ;
 wire \inv_in[2483] ;
 wire \inv_in[2484] ;
 wire \inv_in[2485] ;
 wire \inv_in[2486] ;
 wire \inv_in[2487] ;
 wire \inv_in[2488] ;
 wire \inv_in[2489] ;
 wire \inv_in[248] ;
 wire \inv_in[2490] ;
 wire \inv_in[2491] ;
 wire \inv_in[2492] ;
 wire \inv_in[2493] ;
 wire \inv_in[2494] ;
 wire \inv_in[2495] ;
 wire \inv_in[2496] ;
 wire \inv_in[2497] ;
 wire \inv_in[2498] ;
 wire \inv_in[2499] ;
 wire \inv_in[249] ;
 wire \inv_in[24] ;
 wire \inv_in[2500] ;
 wire \inv_in[2501] ;
 wire \inv_in[2502] ;
 wire \inv_in[2503] ;
 wire \inv_in[2504] ;
 wire \inv_in[2505] ;
 wire \inv_in[2506] ;
 wire \inv_in[2507] ;
 wire \inv_in[2508] ;
 wire \inv_in[2509] ;
 wire \inv_in[250] ;
 wire \inv_in[2510] ;
 wire \inv_in[2511] ;
 wire \inv_in[2512] ;
 wire \inv_in[2513] ;
 wire \inv_in[2514] ;
 wire \inv_in[2515] ;
 wire \inv_in[2516] ;
 wire \inv_in[2517] ;
 wire \inv_in[2518] ;
 wire \inv_in[2519] ;
 wire \inv_in[251] ;
 wire \inv_in[2520] ;
 wire \inv_in[2521] ;
 wire \inv_in[2522] ;
 wire \inv_in[2523] ;
 wire \inv_in[2524] ;
 wire \inv_in[2525] ;
 wire \inv_in[2526] ;
 wire \inv_in[2527] ;
 wire \inv_in[2528] ;
 wire \inv_in[2529] ;
 wire \inv_in[252] ;
 wire \inv_in[2530] ;
 wire \inv_in[2531] ;
 wire \inv_in[2532] ;
 wire \inv_in[2533] ;
 wire \inv_in[2534] ;
 wire \inv_in[2535] ;
 wire \inv_in[2536] ;
 wire \inv_in[2537] ;
 wire \inv_in[2538] ;
 wire \inv_in[2539] ;
 wire \inv_in[253] ;
 wire \inv_in[2540] ;
 wire \inv_in[2541] ;
 wire \inv_in[2542] ;
 wire \inv_in[2543] ;
 wire \inv_in[2544] ;
 wire \inv_in[2545] ;
 wire \inv_in[2546] ;
 wire \inv_in[2547] ;
 wire \inv_in[2548] ;
 wire \inv_in[2549] ;
 wire \inv_in[254] ;
 wire \inv_in[2550] ;
 wire \inv_in[2551] ;
 wire \inv_in[2552] ;
 wire \inv_in[2553] ;
 wire \inv_in[2554] ;
 wire \inv_in[2555] ;
 wire \inv_in[2556] ;
 wire \inv_in[2557] ;
 wire \inv_in[2558] ;
 wire \inv_in[2559] ;
 wire \inv_in[255] ;
 wire \inv_in[2560] ;
 wire \inv_in[2561] ;
 wire \inv_in[2562] ;
 wire \inv_in[2563] ;
 wire \inv_in[2564] ;
 wire \inv_in[2565] ;
 wire \inv_in[2566] ;
 wire \inv_in[2567] ;
 wire \inv_in[2568] ;
 wire \inv_in[2569] ;
 wire \inv_in[256] ;
 wire \inv_in[2570] ;
 wire \inv_in[2571] ;
 wire \inv_in[2572] ;
 wire \inv_in[2573] ;
 wire \inv_in[2574] ;
 wire \inv_in[2575] ;
 wire \inv_in[2576] ;
 wire \inv_in[2577] ;
 wire \inv_in[2578] ;
 wire \inv_in[2579] ;
 wire \inv_in[257] ;
 wire \inv_in[2580] ;
 wire \inv_in[2581] ;
 wire \inv_in[2582] ;
 wire \inv_in[2583] ;
 wire \inv_in[2584] ;
 wire \inv_in[2585] ;
 wire \inv_in[2586] ;
 wire \inv_in[2587] ;
 wire \inv_in[2588] ;
 wire \inv_in[2589] ;
 wire \inv_in[258] ;
 wire \inv_in[2590] ;
 wire \inv_in[2591] ;
 wire \inv_in[2592] ;
 wire \inv_in[2593] ;
 wire \inv_in[2594] ;
 wire \inv_in[2595] ;
 wire \inv_in[2596] ;
 wire \inv_in[2597] ;
 wire \inv_in[2598] ;
 wire \inv_in[2599] ;
 wire \inv_in[259] ;
 wire \inv_in[25] ;
 wire \inv_in[2600] ;
 wire \inv_in[2601] ;
 wire \inv_in[2602] ;
 wire \inv_in[2603] ;
 wire \inv_in[2604] ;
 wire \inv_in[2605] ;
 wire \inv_in[2606] ;
 wire \inv_in[2607] ;
 wire \inv_in[2608] ;
 wire \inv_in[2609] ;
 wire \inv_in[260] ;
 wire \inv_in[2610] ;
 wire \inv_in[2611] ;
 wire \inv_in[2612] ;
 wire \inv_in[2613] ;
 wire \inv_in[2614] ;
 wire \inv_in[2615] ;
 wire \inv_in[2616] ;
 wire \inv_in[2617] ;
 wire \inv_in[2618] ;
 wire \inv_in[2619] ;
 wire \inv_in[261] ;
 wire \inv_in[2620] ;
 wire \inv_in[2621] ;
 wire \inv_in[2622] ;
 wire \inv_in[2623] ;
 wire \inv_in[2624] ;
 wire \inv_in[2625] ;
 wire \inv_in[2626] ;
 wire \inv_in[2627] ;
 wire \inv_in[2628] ;
 wire \inv_in[2629] ;
 wire \inv_in[262] ;
 wire \inv_in[2630] ;
 wire \inv_in[2631] ;
 wire \inv_in[2632] ;
 wire \inv_in[2633] ;
 wire \inv_in[2634] ;
 wire \inv_in[2635] ;
 wire \inv_in[2636] ;
 wire \inv_in[2637] ;
 wire \inv_in[2638] ;
 wire \inv_in[2639] ;
 wire \inv_in[263] ;
 wire \inv_in[2640] ;
 wire \inv_in[2641] ;
 wire \inv_in[2642] ;
 wire \inv_in[2643] ;
 wire \inv_in[2644] ;
 wire \inv_in[2645] ;
 wire \inv_in[2646] ;
 wire \inv_in[2647] ;
 wire \inv_in[2648] ;
 wire \inv_in[2649] ;
 wire \inv_in[264] ;
 wire \inv_in[2650] ;
 wire \inv_in[2651] ;
 wire \inv_in[2652] ;
 wire \inv_in[2653] ;
 wire \inv_in[2654] ;
 wire \inv_in[2655] ;
 wire \inv_in[2656] ;
 wire \inv_in[2657] ;
 wire \inv_in[2658] ;
 wire \inv_in[2659] ;
 wire \inv_in[265] ;
 wire \inv_in[2660] ;
 wire \inv_in[2661] ;
 wire \inv_in[2662] ;
 wire \inv_in[2663] ;
 wire \inv_in[2664] ;
 wire \inv_in[2665] ;
 wire \inv_in[2666] ;
 wire \inv_in[2667] ;
 wire \inv_in[2668] ;
 wire \inv_in[2669] ;
 wire \inv_in[266] ;
 wire \inv_in[2670] ;
 wire \inv_in[2671] ;
 wire \inv_in[2672] ;
 wire \inv_in[2673] ;
 wire \inv_in[2674] ;
 wire \inv_in[2675] ;
 wire \inv_in[2676] ;
 wire \inv_in[2677] ;
 wire \inv_in[2678] ;
 wire \inv_in[2679] ;
 wire \inv_in[267] ;
 wire \inv_in[2680] ;
 wire \inv_in[2681] ;
 wire \inv_in[2682] ;
 wire \inv_in[2683] ;
 wire \inv_in[2684] ;
 wire \inv_in[2685] ;
 wire \inv_in[2686] ;
 wire \inv_in[2687] ;
 wire \inv_in[2688] ;
 wire \inv_in[2689] ;
 wire \inv_in[268] ;
 wire \inv_in[2690] ;
 wire \inv_in[2691] ;
 wire \inv_in[2692] ;
 wire \inv_in[2693] ;
 wire \inv_in[2694] ;
 wire \inv_in[2695] ;
 wire \inv_in[2696] ;
 wire \inv_in[2697] ;
 wire \inv_in[2698] ;
 wire \inv_in[2699] ;
 wire \inv_in[269] ;
 wire \inv_in[26] ;
 wire \inv_in[2700] ;
 wire \inv_in[2701] ;
 wire \inv_in[2702] ;
 wire \inv_in[2703] ;
 wire \inv_in[2704] ;
 wire \inv_in[2705] ;
 wire \inv_in[2706] ;
 wire \inv_in[2707] ;
 wire \inv_in[2708] ;
 wire \inv_in[2709] ;
 wire \inv_in[270] ;
 wire \inv_in[2710] ;
 wire \inv_in[2711] ;
 wire \inv_in[2712] ;
 wire \inv_in[2713] ;
 wire \inv_in[2714] ;
 wire \inv_in[2715] ;
 wire \inv_in[2716] ;
 wire \inv_in[2717] ;
 wire \inv_in[2718] ;
 wire \inv_in[2719] ;
 wire \inv_in[271] ;
 wire \inv_in[2720] ;
 wire \inv_in[2721] ;
 wire \inv_in[2722] ;
 wire \inv_in[2723] ;
 wire \inv_in[2724] ;
 wire \inv_in[2725] ;
 wire \inv_in[2726] ;
 wire \inv_in[2727] ;
 wire \inv_in[2728] ;
 wire \inv_in[2729] ;
 wire \inv_in[272] ;
 wire \inv_in[2730] ;
 wire \inv_in[2731] ;
 wire \inv_in[2732] ;
 wire \inv_in[2733] ;
 wire \inv_in[2734] ;
 wire \inv_in[2735] ;
 wire \inv_in[2736] ;
 wire \inv_in[2737] ;
 wire \inv_in[2738] ;
 wire \inv_in[2739] ;
 wire \inv_in[273] ;
 wire \inv_in[2740] ;
 wire \inv_in[2741] ;
 wire \inv_in[2742] ;
 wire \inv_in[2743] ;
 wire \inv_in[2744] ;
 wire \inv_in[2745] ;
 wire \inv_in[2746] ;
 wire \inv_in[2747] ;
 wire \inv_in[2748] ;
 wire \inv_in[2749] ;
 wire \inv_in[274] ;
 wire \inv_in[2750] ;
 wire \inv_in[2751] ;
 wire \inv_in[2752] ;
 wire \inv_in[2753] ;
 wire \inv_in[2754] ;
 wire \inv_in[2755] ;
 wire \inv_in[2756] ;
 wire \inv_in[2757] ;
 wire \inv_in[2758] ;
 wire \inv_in[2759] ;
 wire \inv_in[275] ;
 wire \inv_in[2760] ;
 wire \inv_in[2761] ;
 wire \inv_in[2762] ;
 wire \inv_in[2763] ;
 wire \inv_in[2764] ;
 wire \inv_in[2765] ;
 wire \inv_in[2766] ;
 wire \inv_in[2767] ;
 wire \inv_in[2768] ;
 wire \inv_in[2769] ;
 wire \inv_in[276] ;
 wire \inv_in[2770] ;
 wire \inv_in[2771] ;
 wire \inv_in[2772] ;
 wire \inv_in[2773] ;
 wire \inv_in[2774] ;
 wire \inv_in[2775] ;
 wire \inv_in[2776] ;
 wire \inv_in[2777] ;
 wire \inv_in[2778] ;
 wire \inv_in[2779] ;
 wire \inv_in[277] ;
 wire \inv_in[2780] ;
 wire \inv_in[2781] ;
 wire \inv_in[2782] ;
 wire \inv_in[2783] ;
 wire \inv_in[2784] ;
 wire \inv_in[2785] ;
 wire \inv_in[2786] ;
 wire \inv_in[2787] ;
 wire \inv_in[2788] ;
 wire \inv_in[2789] ;
 wire \inv_in[278] ;
 wire \inv_in[2790] ;
 wire \inv_in[2791] ;
 wire \inv_in[2792] ;
 wire \inv_in[2793] ;
 wire \inv_in[2794] ;
 wire \inv_in[2795] ;
 wire \inv_in[2796] ;
 wire \inv_in[2797] ;
 wire \inv_in[2798] ;
 wire \inv_in[2799] ;
 wire \inv_in[279] ;
 wire \inv_in[27] ;
 wire \inv_in[2800] ;
 wire \inv_in[2801] ;
 wire \inv_in[2802] ;
 wire \inv_in[2803] ;
 wire \inv_in[2804] ;
 wire \inv_in[2805] ;
 wire \inv_in[2806] ;
 wire \inv_in[2807] ;
 wire \inv_in[2808] ;
 wire \inv_in[2809] ;
 wire \inv_in[280] ;
 wire \inv_in[2810] ;
 wire \inv_in[2811] ;
 wire \inv_in[2812] ;
 wire \inv_in[2813] ;
 wire \inv_in[2814] ;
 wire \inv_in[2815] ;
 wire \inv_in[2816] ;
 wire \inv_in[2817] ;
 wire \inv_in[2818] ;
 wire \inv_in[2819] ;
 wire \inv_in[281] ;
 wire \inv_in[2820] ;
 wire \inv_in[2821] ;
 wire \inv_in[2822] ;
 wire \inv_in[2823] ;
 wire \inv_in[2824] ;
 wire \inv_in[2825] ;
 wire \inv_in[2826] ;
 wire \inv_in[2827] ;
 wire \inv_in[2828] ;
 wire \inv_in[2829] ;
 wire \inv_in[282] ;
 wire \inv_in[2830] ;
 wire \inv_in[2831] ;
 wire \inv_in[2832] ;
 wire \inv_in[2833] ;
 wire \inv_in[2834] ;
 wire \inv_in[2835] ;
 wire \inv_in[2836] ;
 wire \inv_in[2837] ;
 wire \inv_in[2838] ;
 wire \inv_in[2839] ;
 wire \inv_in[283] ;
 wire \inv_in[2840] ;
 wire \inv_in[2841] ;
 wire \inv_in[2842] ;
 wire \inv_in[2843] ;
 wire \inv_in[2844] ;
 wire \inv_in[2845] ;
 wire \inv_in[2846] ;
 wire \inv_in[2847] ;
 wire \inv_in[2848] ;
 wire \inv_in[2849] ;
 wire \inv_in[284] ;
 wire \inv_in[2850] ;
 wire \inv_in[2851] ;
 wire \inv_in[2852] ;
 wire \inv_in[2853] ;
 wire \inv_in[2854] ;
 wire \inv_in[2855] ;
 wire \inv_in[2856] ;
 wire \inv_in[2857] ;
 wire \inv_in[2858] ;
 wire \inv_in[2859] ;
 wire \inv_in[285] ;
 wire \inv_in[2860] ;
 wire \inv_in[2861] ;
 wire \inv_in[2862] ;
 wire \inv_in[2863] ;
 wire \inv_in[2864] ;
 wire \inv_in[2865] ;
 wire \inv_in[2866] ;
 wire \inv_in[2867] ;
 wire \inv_in[2868] ;
 wire \inv_in[2869] ;
 wire \inv_in[286] ;
 wire \inv_in[2870] ;
 wire \inv_in[2871] ;
 wire \inv_in[2872] ;
 wire \inv_in[2873] ;
 wire \inv_in[2874] ;
 wire \inv_in[2875] ;
 wire \inv_in[2876] ;
 wire \inv_in[2877] ;
 wire \inv_in[2878] ;
 wire \inv_in[2879] ;
 wire \inv_in[287] ;
 wire \inv_in[2880] ;
 wire \inv_in[2881] ;
 wire \inv_in[2882] ;
 wire \inv_in[2883] ;
 wire \inv_in[2884] ;
 wire \inv_in[2885] ;
 wire \inv_in[2886] ;
 wire \inv_in[2887] ;
 wire \inv_in[2888] ;
 wire \inv_in[2889] ;
 wire \inv_in[288] ;
 wire \inv_in[2890] ;
 wire \inv_in[2891] ;
 wire \inv_in[2892] ;
 wire \inv_in[2893] ;
 wire \inv_in[2894] ;
 wire \inv_in[2895] ;
 wire \inv_in[2896] ;
 wire \inv_in[2897] ;
 wire \inv_in[2898] ;
 wire \inv_in[2899] ;
 wire \inv_in[289] ;
 wire \inv_in[28] ;
 wire \inv_in[2900] ;
 wire \inv_in[2901] ;
 wire \inv_in[2902] ;
 wire \inv_in[2903] ;
 wire \inv_in[2904] ;
 wire \inv_in[2905] ;
 wire \inv_in[2906] ;
 wire \inv_in[2907] ;
 wire \inv_in[2908] ;
 wire \inv_in[2909] ;
 wire \inv_in[290] ;
 wire \inv_in[2910] ;
 wire \inv_in[2911] ;
 wire \inv_in[2912] ;
 wire \inv_in[2913] ;
 wire \inv_in[2914] ;
 wire \inv_in[2915] ;
 wire \inv_in[2916] ;
 wire \inv_in[2917] ;
 wire \inv_in[2918] ;
 wire \inv_in[2919] ;
 wire \inv_in[291] ;
 wire \inv_in[2920] ;
 wire \inv_in[2921] ;
 wire \inv_in[2922] ;
 wire \inv_in[2923] ;
 wire \inv_in[2924] ;
 wire \inv_in[2925] ;
 wire \inv_in[2926] ;
 wire \inv_in[2927] ;
 wire \inv_in[2928] ;
 wire \inv_in[2929] ;
 wire \inv_in[292] ;
 wire \inv_in[2930] ;
 wire \inv_in[2931] ;
 wire \inv_in[2932] ;
 wire \inv_in[2933] ;
 wire \inv_in[2934] ;
 wire \inv_in[2935] ;
 wire \inv_in[2936] ;
 wire \inv_in[2937] ;
 wire \inv_in[2938] ;
 wire \inv_in[2939] ;
 wire \inv_in[293] ;
 wire \inv_in[2940] ;
 wire \inv_in[2941] ;
 wire \inv_in[2942] ;
 wire \inv_in[2943] ;
 wire \inv_in[2944] ;
 wire \inv_in[2945] ;
 wire \inv_in[2946] ;
 wire \inv_in[2947] ;
 wire \inv_in[2948] ;
 wire \inv_in[2949] ;
 wire \inv_in[294] ;
 wire \inv_in[2950] ;
 wire \inv_in[2951] ;
 wire \inv_in[2952] ;
 wire \inv_in[2953] ;
 wire \inv_in[2954] ;
 wire \inv_in[2955] ;
 wire \inv_in[2956] ;
 wire \inv_in[2957] ;
 wire \inv_in[2958] ;
 wire \inv_in[2959] ;
 wire \inv_in[295] ;
 wire \inv_in[2960] ;
 wire \inv_in[2961] ;
 wire \inv_in[2962] ;
 wire \inv_in[2963] ;
 wire \inv_in[2964] ;
 wire \inv_in[2965] ;
 wire \inv_in[2966] ;
 wire \inv_in[2967] ;
 wire \inv_in[2968] ;
 wire \inv_in[2969] ;
 wire \inv_in[296] ;
 wire \inv_in[2970] ;
 wire \inv_in[2971] ;
 wire \inv_in[2972] ;
 wire \inv_in[2973] ;
 wire \inv_in[2974] ;
 wire \inv_in[2975] ;
 wire \inv_in[2976] ;
 wire \inv_in[2977] ;
 wire \inv_in[2978] ;
 wire \inv_in[2979] ;
 wire \inv_in[297] ;
 wire \inv_in[2980] ;
 wire \inv_in[2981] ;
 wire \inv_in[2982] ;
 wire \inv_in[2983] ;
 wire \inv_in[2984] ;
 wire \inv_in[2985] ;
 wire \inv_in[2986] ;
 wire \inv_in[2987] ;
 wire \inv_in[2988] ;
 wire \inv_in[2989] ;
 wire \inv_in[298] ;
 wire \inv_in[2990] ;
 wire \inv_in[2991] ;
 wire \inv_in[2992] ;
 wire \inv_in[2993] ;
 wire \inv_in[2994] ;
 wire \inv_in[2995] ;
 wire \inv_in[2996] ;
 wire \inv_in[2997] ;
 wire \inv_in[2998] ;
 wire \inv_in[2999] ;
 wire \inv_in[299] ;
 wire \inv_in[29] ;
 wire \inv_in[2] ;
 wire \inv_in[3000] ;
 wire \inv_in[3001] ;
 wire \inv_in[3002] ;
 wire \inv_in[3003] ;
 wire \inv_in[3004] ;
 wire \inv_in[3005] ;
 wire \inv_in[3006] ;
 wire \inv_in[3007] ;
 wire \inv_in[3008] ;
 wire \inv_in[3009] ;
 wire \inv_in[300] ;
 wire \inv_in[3010] ;
 wire \inv_in[3011] ;
 wire \inv_in[3012] ;
 wire \inv_in[3013] ;
 wire \inv_in[3014] ;
 wire \inv_in[3015] ;
 wire \inv_in[3016] ;
 wire \inv_in[3017] ;
 wire \inv_in[3018] ;
 wire \inv_in[3019] ;
 wire \inv_in[301] ;
 wire \inv_in[3020] ;
 wire \inv_in[3021] ;
 wire \inv_in[3022] ;
 wire \inv_in[3023] ;
 wire \inv_in[3024] ;
 wire \inv_in[3025] ;
 wire \inv_in[3026] ;
 wire \inv_in[3027] ;
 wire \inv_in[3028] ;
 wire \inv_in[3029] ;
 wire \inv_in[302] ;
 wire \inv_in[3030] ;
 wire \inv_in[3031] ;
 wire \inv_in[3032] ;
 wire \inv_in[3033] ;
 wire \inv_in[3034] ;
 wire \inv_in[3035] ;
 wire \inv_in[3036] ;
 wire \inv_in[3037] ;
 wire \inv_in[3038] ;
 wire \inv_in[3039] ;
 wire \inv_in[303] ;
 wire \inv_in[3040] ;
 wire \inv_in[3041] ;
 wire \inv_in[3042] ;
 wire \inv_in[3043] ;
 wire \inv_in[3044] ;
 wire \inv_in[3045] ;
 wire \inv_in[3046] ;
 wire \inv_in[3047] ;
 wire \inv_in[3048] ;
 wire \inv_in[3049] ;
 wire \inv_in[304] ;
 wire \inv_in[3050] ;
 wire \inv_in[3051] ;
 wire \inv_in[3052] ;
 wire \inv_in[3053] ;
 wire \inv_in[3054] ;
 wire \inv_in[3055] ;
 wire \inv_in[3056] ;
 wire \inv_in[3057] ;
 wire \inv_in[3058] ;
 wire \inv_in[3059] ;
 wire \inv_in[305] ;
 wire \inv_in[3060] ;
 wire \inv_in[3061] ;
 wire \inv_in[3062] ;
 wire \inv_in[3063] ;
 wire \inv_in[3064] ;
 wire \inv_in[3065] ;
 wire \inv_in[3066] ;
 wire \inv_in[3067] ;
 wire \inv_in[3068] ;
 wire \inv_in[3069] ;
 wire \inv_in[306] ;
 wire \inv_in[3070] ;
 wire \inv_in[3071] ;
 wire \inv_in[3072] ;
 wire \inv_in[3073] ;
 wire \inv_in[3074] ;
 wire \inv_in[3075] ;
 wire \inv_in[3076] ;
 wire \inv_in[3077] ;
 wire \inv_in[3078] ;
 wire \inv_in[3079] ;
 wire \inv_in[307] ;
 wire \inv_in[3080] ;
 wire \inv_in[3081] ;
 wire \inv_in[3082] ;
 wire \inv_in[3083] ;
 wire \inv_in[3084] ;
 wire \inv_in[3085] ;
 wire \inv_in[3086] ;
 wire \inv_in[3087] ;
 wire \inv_in[3088] ;
 wire \inv_in[3089] ;
 wire \inv_in[308] ;
 wire \inv_in[3090] ;
 wire \inv_in[3091] ;
 wire \inv_in[3092] ;
 wire \inv_in[3093] ;
 wire \inv_in[3094] ;
 wire \inv_in[3095] ;
 wire \inv_in[3096] ;
 wire \inv_in[3097] ;
 wire \inv_in[3098] ;
 wire \inv_in[3099] ;
 wire \inv_in[309] ;
 wire \inv_in[30] ;
 wire \inv_in[3100] ;
 wire \inv_in[3101] ;
 wire \inv_in[3102] ;
 wire \inv_in[3103] ;
 wire \inv_in[3104] ;
 wire \inv_in[3105] ;
 wire \inv_in[3106] ;
 wire \inv_in[3107] ;
 wire \inv_in[3108] ;
 wire \inv_in[3109] ;
 wire \inv_in[310] ;
 wire \inv_in[3110] ;
 wire \inv_in[3111] ;
 wire \inv_in[3112] ;
 wire \inv_in[3113] ;
 wire \inv_in[3114] ;
 wire \inv_in[3115] ;
 wire \inv_in[3116] ;
 wire \inv_in[3117] ;
 wire \inv_in[3118] ;
 wire \inv_in[3119] ;
 wire \inv_in[311] ;
 wire \inv_in[3120] ;
 wire \inv_in[3121] ;
 wire \inv_in[3122] ;
 wire \inv_in[3123] ;
 wire \inv_in[3124] ;
 wire \inv_in[3125] ;
 wire \inv_in[3126] ;
 wire \inv_in[3127] ;
 wire \inv_in[3128] ;
 wire \inv_in[3129] ;
 wire \inv_in[312] ;
 wire \inv_in[3130] ;
 wire \inv_in[3131] ;
 wire \inv_in[3132] ;
 wire \inv_in[3133] ;
 wire \inv_in[3134] ;
 wire \inv_in[3135] ;
 wire \inv_in[3136] ;
 wire \inv_in[3137] ;
 wire \inv_in[3138] ;
 wire \inv_in[3139] ;
 wire \inv_in[313] ;
 wire \inv_in[3140] ;
 wire \inv_in[3141] ;
 wire \inv_in[3142] ;
 wire \inv_in[3143] ;
 wire \inv_in[3144] ;
 wire \inv_in[3145] ;
 wire \inv_in[3146] ;
 wire \inv_in[3147] ;
 wire \inv_in[3148] ;
 wire \inv_in[3149] ;
 wire \inv_in[314] ;
 wire \inv_in[3150] ;
 wire \inv_in[3151] ;
 wire \inv_in[3152] ;
 wire \inv_in[3153] ;
 wire \inv_in[3154] ;
 wire \inv_in[3155] ;
 wire \inv_in[3156] ;
 wire \inv_in[3157] ;
 wire \inv_in[3158] ;
 wire \inv_in[3159] ;
 wire \inv_in[315] ;
 wire \inv_in[3160] ;
 wire \inv_in[3161] ;
 wire \inv_in[3162] ;
 wire \inv_in[3163] ;
 wire \inv_in[3164] ;
 wire \inv_in[3165] ;
 wire \inv_in[3166] ;
 wire \inv_in[3167] ;
 wire \inv_in[3168] ;
 wire \inv_in[3169] ;
 wire \inv_in[316] ;
 wire \inv_in[3170] ;
 wire \inv_in[3171] ;
 wire \inv_in[3172] ;
 wire \inv_in[3173] ;
 wire \inv_in[3174] ;
 wire \inv_in[3175] ;
 wire \inv_in[3176] ;
 wire \inv_in[3177] ;
 wire \inv_in[3178] ;
 wire \inv_in[3179] ;
 wire \inv_in[317] ;
 wire \inv_in[3180] ;
 wire \inv_in[3181] ;
 wire \inv_in[3182] ;
 wire \inv_in[3183] ;
 wire \inv_in[3184] ;
 wire \inv_in[3185] ;
 wire \inv_in[3186] ;
 wire \inv_in[3187] ;
 wire \inv_in[3188] ;
 wire \inv_in[3189] ;
 wire \inv_in[318] ;
 wire \inv_in[3190] ;
 wire \inv_in[3191] ;
 wire \inv_in[3192] ;
 wire \inv_in[3193] ;
 wire \inv_in[3194] ;
 wire \inv_in[3195] ;
 wire \inv_in[3196] ;
 wire \inv_in[3197] ;
 wire \inv_in[3198] ;
 wire \inv_in[3199] ;
 wire \inv_in[319] ;
 wire \inv_in[31] ;
 wire \inv_in[3200] ;
 wire \inv_in[3201] ;
 wire \inv_in[3202] ;
 wire \inv_in[3203] ;
 wire \inv_in[3204] ;
 wire \inv_in[3205] ;
 wire \inv_in[3206] ;
 wire \inv_in[3207] ;
 wire \inv_in[3208] ;
 wire \inv_in[3209] ;
 wire \inv_in[320] ;
 wire \inv_in[3210] ;
 wire \inv_in[3211] ;
 wire \inv_in[3212] ;
 wire \inv_in[3213] ;
 wire \inv_in[3214] ;
 wire \inv_in[3215] ;
 wire \inv_in[3216] ;
 wire \inv_in[3217] ;
 wire \inv_in[3218] ;
 wire \inv_in[3219] ;
 wire \inv_in[321] ;
 wire \inv_in[3220] ;
 wire \inv_in[3221] ;
 wire \inv_in[3222] ;
 wire \inv_in[3223] ;
 wire \inv_in[3224] ;
 wire \inv_in[3225] ;
 wire \inv_in[3226] ;
 wire \inv_in[3227] ;
 wire \inv_in[3228] ;
 wire \inv_in[3229] ;
 wire \inv_in[322] ;
 wire \inv_in[3230] ;
 wire \inv_in[3231] ;
 wire \inv_in[3232] ;
 wire \inv_in[3233] ;
 wire \inv_in[3234] ;
 wire \inv_in[3235] ;
 wire \inv_in[3236] ;
 wire \inv_in[3237] ;
 wire \inv_in[3238] ;
 wire \inv_in[3239] ;
 wire \inv_in[323] ;
 wire \inv_in[3240] ;
 wire \inv_in[3241] ;
 wire \inv_in[3242] ;
 wire \inv_in[3243] ;
 wire \inv_in[3244] ;
 wire \inv_in[3245] ;
 wire \inv_in[3246] ;
 wire \inv_in[3247] ;
 wire \inv_in[3248] ;
 wire \inv_in[3249] ;
 wire \inv_in[324] ;
 wire \inv_in[3250] ;
 wire \inv_in[3251] ;
 wire \inv_in[3252] ;
 wire \inv_in[3253] ;
 wire \inv_in[3254] ;
 wire \inv_in[3255] ;
 wire \inv_in[3256] ;
 wire \inv_in[3257] ;
 wire \inv_in[3258] ;
 wire \inv_in[3259] ;
 wire \inv_in[325] ;
 wire \inv_in[3260] ;
 wire \inv_in[3261] ;
 wire \inv_in[3262] ;
 wire \inv_in[3263] ;
 wire \inv_in[3264] ;
 wire \inv_in[3265] ;
 wire \inv_in[3266] ;
 wire \inv_in[3267] ;
 wire \inv_in[3268] ;
 wire \inv_in[3269] ;
 wire \inv_in[326] ;
 wire \inv_in[3270] ;
 wire \inv_in[3271] ;
 wire \inv_in[3272] ;
 wire \inv_in[3273] ;
 wire \inv_in[3274] ;
 wire \inv_in[3275] ;
 wire \inv_in[3276] ;
 wire \inv_in[3277] ;
 wire \inv_in[3278] ;
 wire \inv_in[3279] ;
 wire \inv_in[327] ;
 wire \inv_in[3280] ;
 wire \inv_in[3281] ;
 wire \inv_in[3282] ;
 wire \inv_in[3283] ;
 wire \inv_in[3284] ;
 wire \inv_in[3285] ;
 wire \inv_in[3286] ;
 wire \inv_in[3287] ;
 wire \inv_in[3288] ;
 wire \inv_in[3289] ;
 wire \inv_in[328] ;
 wire \inv_in[3290] ;
 wire \inv_in[3291] ;
 wire \inv_in[3292] ;
 wire \inv_in[3293] ;
 wire \inv_in[3294] ;
 wire \inv_in[3295] ;
 wire \inv_in[3296] ;
 wire \inv_in[3297] ;
 wire \inv_in[3298] ;
 wire \inv_in[3299] ;
 wire \inv_in[329] ;
 wire \inv_in[32] ;
 wire \inv_in[3300] ;
 wire \inv_in[3301] ;
 wire \inv_in[3302] ;
 wire \inv_in[3303] ;
 wire \inv_in[3304] ;
 wire \inv_in[3305] ;
 wire \inv_in[3306] ;
 wire \inv_in[3307] ;
 wire \inv_in[3308] ;
 wire \inv_in[3309] ;
 wire \inv_in[330] ;
 wire \inv_in[3310] ;
 wire \inv_in[3311] ;
 wire \inv_in[3312] ;
 wire \inv_in[3313] ;
 wire \inv_in[3314] ;
 wire \inv_in[3315] ;
 wire \inv_in[3316] ;
 wire \inv_in[3317] ;
 wire \inv_in[3318] ;
 wire \inv_in[3319] ;
 wire \inv_in[331] ;
 wire \inv_in[3320] ;
 wire \inv_in[3321] ;
 wire \inv_in[3322] ;
 wire \inv_in[3323] ;
 wire \inv_in[3324] ;
 wire \inv_in[3325] ;
 wire \inv_in[3326] ;
 wire \inv_in[3327] ;
 wire \inv_in[3328] ;
 wire \inv_in[3329] ;
 wire \inv_in[332] ;
 wire \inv_in[3330] ;
 wire \inv_in[3331] ;
 wire \inv_in[3332] ;
 wire \inv_in[3333] ;
 wire \inv_in[3334] ;
 wire \inv_in[3335] ;
 wire \inv_in[3336] ;
 wire \inv_in[3337] ;
 wire \inv_in[3338] ;
 wire \inv_in[3339] ;
 wire \inv_in[333] ;
 wire \inv_in[3340] ;
 wire \inv_in[3341] ;
 wire \inv_in[3342] ;
 wire \inv_in[3343] ;
 wire \inv_in[3344] ;
 wire \inv_in[3345] ;
 wire \inv_in[3346] ;
 wire \inv_in[3347] ;
 wire \inv_in[3348] ;
 wire \inv_in[3349] ;
 wire \inv_in[334] ;
 wire \inv_in[3350] ;
 wire \inv_in[3351] ;
 wire \inv_in[3352] ;
 wire \inv_in[3353] ;
 wire \inv_in[3354] ;
 wire \inv_in[3355] ;
 wire \inv_in[3356] ;
 wire \inv_in[3357] ;
 wire \inv_in[3358] ;
 wire \inv_in[3359] ;
 wire \inv_in[335] ;
 wire \inv_in[3360] ;
 wire \inv_in[3361] ;
 wire \inv_in[3362] ;
 wire \inv_in[3363] ;
 wire \inv_in[3364] ;
 wire \inv_in[3365] ;
 wire \inv_in[3366] ;
 wire \inv_in[3367] ;
 wire \inv_in[3368] ;
 wire \inv_in[3369] ;
 wire \inv_in[336] ;
 wire \inv_in[3370] ;
 wire \inv_in[3371] ;
 wire \inv_in[3372] ;
 wire \inv_in[3373] ;
 wire \inv_in[3374] ;
 wire \inv_in[3375] ;
 wire \inv_in[3376] ;
 wire \inv_in[3377] ;
 wire \inv_in[3378] ;
 wire \inv_in[3379] ;
 wire \inv_in[337] ;
 wire \inv_in[3380] ;
 wire \inv_in[3381] ;
 wire \inv_in[3382] ;
 wire \inv_in[3383] ;
 wire \inv_in[3384] ;
 wire \inv_in[3385] ;
 wire \inv_in[3386] ;
 wire \inv_in[3387] ;
 wire \inv_in[3388] ;
 wire \inv_in[3389] ;
 wire \inv_in[338] ;
 wire \inv_in[3390] ;
 wire \inv_in[3391] ;
 wire \inv_in[3392] ;
 wire \inv_in[3393] ;
 wire \inv_in[3394] ;
 wire \inv_in[3395] ;
 wire \inv_in[3396] ;
 wire \inv_in[3397] ;
 wire \inv_in[3398] ;
 wire \inv_in[3399] ;
 wire \inv_in[339] ;
 wire \inv_in[33] ;
 wire \inv_in[3400] ;
 wire \inv_in[3401] ;
 wire \inv_in[3402] ;
 wire \inv_in[3403] ;
 wire \inv_in[3404] ;
 wire \inv_in[3405] ;
 wire \inv_in[3406] ;
 wire \inv_in[3407] ;
 wire \inv_in[3408] ;
 wire \inv_in[3409] ;
 wire \inv_in[340] ;
 wire \inv_in[3410] ;
 wire \inv_in[3411] ;
 wire \inv_in[3412] ;
 wire \inv_in[3413] ;
 wire \inv_in[3414] ;
 wire \inv_in[3415] ;
 wire \inv_in[3416] ;
 wire \inv_in[3417] ;
 wire \inv_in[3418] ;
 wire \inv_in[3419] ;
 wire \inv_in[341] ;
 wire \inv_in[3420] ;
 wire \inv_in[3421] ;
 wire \inv_in[3422] ;
 wire \inv_in[3423] ;
 wire \inv_in[3424] ;
 wire \inv_in[3425] ;
 wire \inv_in[3426] ;
 wire \inv_in[3427] ;
 wire \inv_in[3428] ;
 wire \inv_in[3429] ;
 wire \inv_in[342] ;
 wire \inv_in[3430] ;
 wire \inv_in[3431] ;
 wire \inv_in[3432] ;
 wire \inv_in[3433] ;
 wire \inv_in[3434] ;
 wire \inv_in[3435] ;
 wire \inv_in[3436] ;
 wire \inv_in[3437] ;
 wire \inv_in[3438] ;
 wire \inv_in[3439] ;
 wire \inv_in[343] ;
 wire \inv_in[3440] ;
 wire \inv_in[3441] ;
 wire \inv_in[3442] ;
 wire \inv_in[3443] ;
 wire \inv_in[3444] ;
 wire \inv_in[3445] ;
 wire \inv_in[3446] ;
 wire \inv_in[3447] ;
 wire \inv_in[3448] ;
 wire \inv_in[3449] ;
 wire \inv_in[344] ;
 wire \inv_in[3450] ;
 wire \inv_in[3451] ;
 wire \inv_in[3452] ;
 wire \inv_in[3453] ;
 wire \inv_in[3454] ;
 wire \inv_in[3455] ;
 wire \inv_in[3456] ;
 wire \inv_in[3457] ;
 wire \inv_in[3458] ;
 wire \inv_in[3459] ;
 wire \inv_in[345] ;
 wire \inv_in[3460] ;
 wire \inv_in[3461] ;
 wire \inv_in[3462] ;
 wire \inv_in[3463] ;
 wire \inv_in[3464] ;
 wire \inv_in[3465] ;
 wire \inv_in[3466] ;
 wire \inv_in[3467] ;
 wire \inv_in[3468] ;
 wire \inv_in[3469] ;
 wire \inv_in[346] ;
 wire \inv_in[3470] ;
 wire \inv_in[3471] ;
 wire \inv_in[3472] ;
 wire \inv_in[3473] ;
 wire \inv_in[3474] ;
 wire \inv_in[3475] ;
 wire \inv_in[3476] ;
 wire \inv_in[3477] ;
 wire \inv_in[3478] ;
 wire \inv_in[3479] ;
 wire \inv_in[347] ;
 wire \inv_in[3480] ;
 wire \inv_in[3481] ;
 wire \inv_in[3482] ;
 wire \inv_in[3483] ;
 wire \inv_in[3484] ;
 wire \inv_in[3485] ;
 wire \inv_in[3486] ;
 wire \inv_in[3487] ;
 wire \inv_in[3488] ;
 wire \inv_in[3489] ;
 wire \inv_in[348] ;
 wire \inv_in[3490] ;
 wire \inv_in[3491] ;
 wire \inv_in[3492] ;
 wire \inv_in[3493] ;
 wire \inv_in[3494] ;
 wire \inv_in[3495] ;
 wire \inv_in[3496] ;
 wire \inv_in[3497] ;
 wire \inv_in[3498] ;
 wire \inv_in[3499] ;
 wire \inv_in[349] ;
 wire \inv_in[34] ;
 wire \inv_in[3500] ;
 wire \inv_in[3501] ;
 wire \inv_in[3502] ;
 wire \inv_in[3503] ;
 wire \inv_in[3504] ;
 wire \inv_in[3505] ;
 wire \inv_in[3506] ;
 wire \inv_in[3507] ;
 wire \inv_in[3508] ;
 wire \inv_in[3509] ;
 wire \inv_in[350] ;
 wire \inv_in[3510] ;
 wire \inv_in[3511] ;
 wire \inv_in[3512] ;
 wire \inv_in[3513] ;
 wire \inv_in[3514] ;
 wire \inv_in[3515] ;
 wire \inv_in[3516] ;
 wire \inv_in[3517] ;
 wire \inv_in[3518] ;
 wire \inv_in[3519] ;
 wire \inv_in[351] ;
 wire \inv_in[3520] ;
 wire \inv_in[3521] ;
 wire \inv_in[3522] ;
 wire \inv_in[3523] ;
 wire \inv_in[3524] ;
 wire \inv_in[3525] ;
 wire \inv_in[3526] ;
 wire \inv_in[3527] ;
 wire \inv_in[3528] ;
 wire \inv_in[3529] ;
 wire \inv_in[352] ;
 wire \inv_in[3530] ;
 wire \inv_in[3531] ;
 wire \inv_in[3532] ;
 wire \inv_in[3533] ;
 wire \inv_in[3534] ;
 wire \inv_in[3535] ;
 wire \inv_in[3536] ;
 wire \inv_in[3537] ;
 wire \inv_in[3538] ;
 wire \inv_in[3539] ;
 wire \inv_in[353] ;
 wire \inv_in[3540] ;
 wire \inv_in[3541] ;
 wire \inv_in[3542] ;
 wire \inv_in[3543] ;
 wire \inv_in[3544] ;
 wire \inv_in[3545] ;
 wire \inv_in[3546] ;
 wire \inv_in[3547] ;
 wire \inv_in[3548] ;
 wire \inv_in[3549] ;
 wire \inv_in[354] ;
 wire \inv_in[3550] ;
 wire \inv_in[3551] ;
 wire \inv_in[3552] ;
 wire \inv_in[3553] ;
 wire \inv_in[3554] ;
 wire \inv_in[3555] ;
 wire \inv_in[3556] ;
 wire \inv_in[3557] ;
 wire \inv_in[3558] ;
 wire \inv_in[3559] ;
 wire \inv_in[355] ;
 wire \inv_in[3560] ;
 wire \inv_in[3561] ;
 wire \inv_in[3562] ;
 wire \inv_in[3563] ;
 wire \inv_in[3564] ;
 wire \inv_in[3565] ;
 wire \inv_in[3566] ;
 wire \inv_in[3567] ;
 wire \inv_in[3568] ;
 wire \inv_in[3569] ;
 wire \inv_in[356] ;
 wire \inv_in[3570] ;
 wire \inv_in[3571] ;
 wire \inv_in[3572] ;
 wire \inv_in[3573] ;
 wire \inv_in[3574] ;
 wire \inv_in[3575] ;
 wire \inv_in[3576] ;
 wire \inv_in[3577] ;
 wire \inv_in[3578] ;
 wire \inv_in[3579] ;
 wire \inv_in[357] ;
 wire \inv_in[3580] ;
 wire \inv_in[3581] ;
 wire \inv_in[3582] ;
 wire \inv_in[3583] ;
 wire \inv_in[3584] ;
 wire \inv_in[3585] ;
 wire \inv_in[3586] ;
 wire \inv_in[3587] ;
 wire \inv_in[3588] ;
 wire \inv_in[3589] ;
 wire \inv_in[358] ;
 wire \inv_in[3590] ;
 wire \inv_in[3591] ;
 wire \inv_in[3592] ;
 wire \inv_in[3593] ;
 wire \inv_in[3594] ;
 wire \inv_in[3595] ;
 wire \inv_in[3596] ;
 wire \inv_in[3597] ;
 wire \inv_in[3598] ;
 wire \inv_in[3599] ;
 wire \inv_in[359] ;
 wire \inv_in[35] ;
 wire \inv_in[3600] ;
 wire \inv_in[3601] ;
 wire \inv_in[3602] ;
 wire \inv_in[3603] ;
 wire \inv_in[3604] ;
 wire \inv_in[3605] ;
 wire \inv_in[3606] ;
 wire \inv_in[3607] ;
 wire \inv_in[3608] ;
 wire \inv_in[3609] ;
 wire \inv_in[360] ;
 wire \inv_in[3610] ;
 wire \inv_in[3611] ;
 wire \inv_in[3612] ;
 wire \inv_in[3613] ;
 wire \inv_in[3614] ;
 wire \inv_in[3615] ;
 wire \inv_in[3616] ;
 wire \inv_in[3617] ;
 wire \inv_in[3618] ;
 wire \inv_in[3619] ;
 wire \inv_in[361] ;
 wire \inv_in[3620] ;
 wire \inv_in[3621] ;
 wire \inv_in[3622] ;
 wire \inv_in[3623] ;
 wire \inv_in[3624] ;
 wire \inv_in[3625] ;
 wire \inv_in[3626] ;
 wire \inv_in[3627] ;
 wire \inv_in[3628] ;
 wire \inv_in[3629] ;
 wire \inv_in[362] ;
 wire \inv_in[3630] ;
 wire \inv_in[3631] ;
 wire \inv_in[3632] ;
 wire \inv_in[3633] ;
 wire \inv_in[3634] ;
 wire \inv_in[3635] ;
 wire \inv_in[3636] ;
 wire \inv_in[3637] ;
 wire \inv_in[3638] ;
 wire \inv_in[3639] ;
 wire \inv_in[363] ;
 wire \inv_in[3640] ;
 wire \inv_in[3641] ;
 wire \inv_in[3642] ;
 wire \inv_in[3643] ;
 wire \inv_in[3644] ;
 wire \inv_in[3645] ;
 wire \inv_in[3646] ;
 wire \inv_in[3647] ;
 wire \inv_in[3648] ;
 wire \inv_in[3649] ;
 wire \inv_in[364] ;
 wire \inv_in[3650] ;
 wire \inv_in[3651] ;
 wire \inv_in[3652] ;
 wire \inv_in[3653] ;
 wire \inv_in[3654] ;
 wire \inv_in[3655] ;
 wire \inv_in[3656] ;
 wire \inv_in[3657] ;
 wire \inv_in[3658] ;
 wire \inv_in[3659] ;
 wire \inv_in[365] ;
 wire \inv_in[3660] ;
 wire \inv_in[3661] ;
 wire \inv_in[3662] ;
 wire \inv_in[3663] ;
 wire \inv_in[3664] ;
 wire \inv_in[3665] ;
 wire \inv_in[3666] ;
 wire \inv_in[3667] ;
 wire \inv_in[3668] ;
 wire \inv_in[3669] ;
 wire \inv_in[366] ;
 wire \inv_in[3670] ;
 wire \inv_in[3671] ;
 wire \inv_in[3672] ;
 wire \inv_in[3673] ;
 wire \inv_in[3674] ;
 wire \inv_in[3675] ;
 wire \inv_in[3676] ;
 wire \inv_in[3677] ;
 wire \inv_in[3678] ;
 wire \inv_in[3679] ;
 wire \inv_in[367] ;
 wire \inv_in[3680] ;
 wire \inv_in[3681] ;
 wire \inv_in[3682] ;
 wire \inv_in[3683] ;
 wire \inv_in[3684] ;
 wire \inv_in[3685] ;
 wire \inv_in[3686] ;
 wire \inv_in[3687] ;
 wire \inv_in[3688] ;
 wire \inv_in[3689] ;
 wire \inv_in[368] ;
 wire \inv_in[3690] ;
 wire \inv_in[3691] ;
 wire \inv_in[3692] ;
 wire \inv_in[3693] ;
 wire \inv_in[3694] ;
 wire \inv_in[3695] ;
 wire \inv_in[3696] ;
 wire \inv_in[3697] ;
 wire \inv_in[3698] ;
 wire \inv_in[3699] ;
 wire \inv_in[369] ;
 wire \inv_in[36] ;
 wire \inv_in[3700] ;
 wire \inv_in[3701] ;
 wire \inv_in[3702] ;
 wire \inv_in[3703] ;
 wire \inv_in[3704] ;
 wire \inv_in[3705] ;
 wire \inv_in[3706] ;
 wire \inv_in[3707] ;
 wire \inv_in[3708] ;
 wire \inv_in[3709] ;
 wire \inv_in[370] ;
 wire \inv_in[3710] ;
 wire \inv_in[3711] ;
 wire \inv_in[3712] ;
 wire \inv_in[3713] ;
 wire \inv_in[3714] ;
 wire \inv_in[3715] ;
 wire \inv_in[3716] ;
 wire \inv_in[3717] ;
 wire \inv_in[3718] ;
 wire \inv_in[3719] ;
 wire \inv_in[371] ;
 wire \inv_in[3720] ;
 wire \inv_in[3721] ;
 wire \inv_in[3722] ;
 wire \inv_in[3723] ;
 wire \inv_in[3724] ;
 wire \inv_in[3725] ;
 wire \inv_in[3726] ;
 wire \inv_in[3727] ;
 wire \inv_in[3728] ;
 wire \inv_in[3729] ;
 wire \inv_in[372] ;
 wire \inv_in[3730] ;
 wire \inv_in[3731] ;
 wire \inv_in[3732] ;
 wire \inv_in[3733] ;
 wire \inv_in[3734] ;
 wire \inv_in[3735] ;
 wire \inv_in[3736] ;
 wire \inv_in[3737] ;
 wire \inv_in[3738] ;
 wire \inv_in[3739] ;
 wire \inv_in[373] ;
 wire \inv_in[3740] ;
 wire \inv_in[3741] ;
 wire \inv_in[3742] ;
 wire \inv_in[3743] ;
 wire \inv_in[3744] ;
 wire \inv_in[3745] ;
 wire \inv_in[3746] ;
 wire \inv_in[3747] ;
 wire \inv_in[3748] ;
 wire \inv_in[3749] ;
 wire \inv_in[374] ;
 wire \inv_in[3750] ;
 wire \inv_in[3751] ;
 wire \inv_in[3752] ;
 wire \inv_in[3753] ;
 wire \inv_in[3754] ;
 wire \inv_in[3755] ;
 wire \inv_in[3756] ;
 wire \inv_in[3757] ;
 wire \inv_in[3758] ;
 wire \inv_in[3759] ;
 wire \inv_in[375] ;
 wire \inv_in[3760] ;
 wire \inv_in[3761] ;
 wire \inv_in[3762] ;
 wire \inv_in[3763] ;
 wire \inv_in[3764] ;
 wire \inv_in[3765] ;
 wire \inv_in[3766] ;
 wire \inv_in[3767] ;
 wire \inv_in[3768] ;
 wire \inv_in[3769] ;
 wire \inv_in[376] ;
 wire \inv_in[3770] ;
 wire \inv_in[3771] ;
 wire \inv_in[3772] ;
 wire \inv_in[3773] ;
 wire \inv_in[3774] ;
 wire \inv_in[3775] ;
 wire \inv_in[3776] ;
 wire \inv_in[3777] ;
 wire \inv_in[3778] ;
 wire \inv_in[3779] ;
 wire \inv_in[377] ;
 wire \inv_in[3780] ;
 wire \inv_in[3781] ;
 wire \inv_in[3782] ;
 wire \inv_in[3783] ;
 wire \inv_in[3784] ;
 wire \inv_in[3785] ;
 wire \inv_in[3786] ;
 wire \inv_in[3787] ;
 wire \inv_in[3788] ;
 wire \inv_in[3789] ;
 wire \inv_in[378] ;
 wire \inv_in[3790] ;
 wire \inv_in[3791] ;
 wire \inv_in[3792] ;
 wire \inv_in[3793] ;
 wire \inv_in[3794] ;
 wire \inv_in[3795] ;
 wire \inv_in[3796] ;
 wire \inv_in[3797] ;
 wire \inv_in[3798] ;
 wire \inv_in[3799] ;
 wire \inv_in[379] ;
 wire \inv_in[37] ;
 wire \inv_in[3800] ;
 wire \inv_in[3801] ;
 wire \inv_in[3802] ;
 wire \inv_in[3803] ;
 wire \inv_in[3804] ;
 wire \inv_in[3805] ;
 wire \inv_in[3806] ;
 wire \inv_in[3807] ;
 wire \inv_in[3808] ;
 wire \inv_in[3809] ;
 wire \inv_in[380] ;
 wire \inv_in[3810] ;
 wire \inv_in[3811] ;
 wire \inv_in[3812] ;
 wire \inv_in[3813] ;
 wire \inv_in[3814] ;
 wire \inv_in[3815] ;
 wire \inv_in[3816] ;
 wire \inv_in[3817] ;
 wire \inv_in[3818] ;
 wire \inv_in[3819] ;
 wire \inv_in[381] ;
 wire \inv_in[3820] ;
 wire \inv_in[3821] ;
 wire \inv_in[3822] ;
 wire \inv_in[3823] ;
 wire \inv_in[3824] ;
 wire \inv_in[3825] ;
 wire \inv_in[3826] ;
 wire \inv_in[3827] ;
 wire \inv_in[3828] ;
 wire \inv_in[3829] ;
 wire \inv_in[382] ;
 wire \inv_in[3830] ;
 wire \inv_in[3831] ;
 wire \inv_in[3832] ;
 wire \inv_in[3833] ;
 wire \inv_in[3834] ;
 wire \inv_in[3835] ;
 wire \inv_in[3836] ;
 wire \inv_in[3837] ;
 wire \inv_in[3838] ;
 wire \inv_in[3839] ;
 wire \inv_in[383] ;
 wire \inv_in[3840] ;
 wire \inv_in[3841] ;
 wire \inv_in[3842] ;
 wire \inv_in[3843] ;
 wire \inv_in[3844] ;
 wire \inv_in[3845] ;
 wire \inv_in[3846] ;
 wire \inv_in[3847] ;
 wire \inv_in[3848] ;
 wire \inv_in[3849] ;
 wire \inv_in[384] ;
 wire \inv_in[3850] ;
 wire \inv_in[3851] ;
 wire \inv_in[3852] ;
 wire \inv_in[385] ;
 wire \inv_in[386] ;
 wire \inv_in[387] ;
 wire \inv_in[388] ;
 wire \inv_in[389] ;
 wire \inv_in[38] ;
 wire \inv_in[390] ;
 wire \inv_in[391] ;
 wire \inv_in[392] ;
 wire \inv_in[393] ;
 wire \inv_in[394] ;
 wire \inv_in[395] ;
 wire \inv_in[396] ;
 wire \inv_in[397] ;
 wire \inv_in[398] ;
 wire \inv_in[399] ;
 wire \inv_in[39] ;
 wire \inv_in[3] ;
 wire \inv_in[400] ;
 wire \inv_in[401] ;
 wire \inv_in[402] ;
 wire \inv_in[403] ;
 wire \inv_in[404] ;
 wire \inv_in[405] ;
 wire \inv_in[406] ;
 wire \inv_in[407] ;
 wire \inv_in[408] ;
 wire \inv_in[409] ;
 wire \inv_in[40] ;
 wire \inv_in[410] ;
 wire \inv_in[411] ;
 wire \inv_in[412] ;
 wire \inv_in[413] ;
 wire \inv_in[414] ;
 wire \inv_in[415] ;
 wire \inv_in[416] ;
 wire \inv_in[417] ;
 wire \inv_in[418] ;
 wire \inv_in[419] ;
 wire \inv_in[41] ;
 wire \inv_in[420] ;
 wire \inv_in[421] ;
 wire \inv_in[422] ;
 wire \inv_in[423] ;
 wire \inv_in[424] ;
 wire \inv_in[425] ;
 wire \inv_in[426] ;
 wire \inv_in[427] ;
 wire \inv_in[428] ;
 wire \inv_in[429] ;
 wire \inv_in[42] ;
 wire \inv_in[430] ;
 wire \inv_in[431] ;
 wire \inv_in[432] ;
 wire \inv_in[433] ;
 wire \inv_in[434] ;
 wire \inv_in[435] ;
 wire \inv_in[436] ;
 wire \inv_in[437] ;
 wire \inv_in[438] ;
 wire \inv_in[439] ;
 wire \inv_in[43] ;
 wire \inv_in[440] ;
 wire \inv_in[441] ;
 wire \inv_in[442] ;
 wire \inv_in[443] ;
 wire \inv_in[444] ;
 wire \inv_in[445] ;
 wire \inv_in[446] ;
 wire \inv_in[447] ;
 wire \inv_in[448] ;
 wire \inv_in[449] ;
 wire \inv_in[44] ;
 wire \inv_in[450] ;
 wire \inv_in[451] ;
 wire \inv_in[452] ;
 wire \inv_in[453] ;
 wire \inv_in[454] ;
 wire \inv_in[455] ;
 wire \inv_in[456] ;
 wire \inv_in[457] ;
 wire \inv_in[458] ;
 wire \inv_in[459] ;
 wire \inv_in[45] ;
 wire \inv_in[460] ;
 wire \inv_in[461] ;
 wire \inv_in[462] ;
 wire \inv_in[463] ;
 wire \inv_in[464] ;
 wire \inv_in[465] ;
 wire \inv_in[466] ;
 wire \inv_in[467] ;
 wire \inv_in[468] ;
 wire \inv_in[469] ;
 wire \inv_in[46] ;
 wire \inv_in[470] ;
 wire \inv_in[471] ;
 wire \inv_in[472] ;
 wire \inv_in[473] ;
 wire \inv_in[474] ;
 wire \inv_in[475] ;
 wire \inv_in[476] ;
 wire \inv_in[477] ;
 wire \inv_in[478] ;
 wire \inv_in[479] ;
 wire \inv_in[47] ;
 wire \inv_in[480] ;
 wire \inv_in[481] ;
 wire \inv_in[482] ;
 wire \inv_in[483] ;
 wire \inv_in[484] ;
 wire \inv_in[485] ;
 wire \inv_in[486] ;
 wire \inv_in[487] ;
 wire \inv_in[488] ;
 wire \inv_in[489] ;
 wire \inv_in[48] ;
 wire \inv_in[490] ;
 wire \inv_in[491] ;
 wire \inv_in[492] ;
 wire \inv_in[493] ;
 wire \inv_in[494] ;
 wire \inv_in[495] ;
 wire \inv_in[496] ;
 wire \inv_in[497] ;
 wire \inv_in[498] ;
 wire \inv_in[499] ;
 wire \inv_in[49] ;
 wire \inv_in[4] ;
 wire \inv_in[500] ;
 wire \inv_in[501] ;
 wire \inv_in[502] ;
 wire \inv_in[503] ;
 wire \inv_in[504] ;
 wire \inv_in[505] ;
 wire \inv_in[506] ;
 wire \inv_in[507] ;
 wire \inv_in[508] ;
 wire \inv_in[509] ;
 wire \inv_in[50] ;
 wire \inv_in[510] ;
 wire \inv_in[511] ;
 wire \inv_in[512] ;
 wire \inv_in[513] ;
 wire \inv_in[514] ;
 wire \inv_in[515] ;
 wire \inv_in[516] ;
 wire \inv_in[517] ;
 wire \inv_in[518] ;
 wire \inv_in[519] ;
 wire \inv_in[51] ;
 wire \inv_in[520] ;
 wire \inv_in[521] ;
 wire \inv_in[522] ;
 wire \inv_in[523] ;
 wire \inv_in[524] ;
 wire \inv_in[525] ;
 wire \inv_in[526] ;
 wire \inv_in[527] ;
 wire \inv_in[528] ;
 wire \inv_in[529] ;
 wire \inv_in[52] ;
 wire \inv_in[530] ;
 wire \inv_in[531] ;
 wire \inv_in[532] ;
 wire \inv_in[533] ;
 wire \inv_in[534] ;
 wire \inv_in[535] ;
 wire \inv_in[536] ;
 wire \inv_in[537] ;
 wire \inv_in[538] ;
 wire \inv_in[539] ;
 wire \inv_in[53] ;
 wire \inv_in[540] ;
 wire \inv_in[541] ;
 wire \inv_in[542] ;
 wire \inv_in[543] ;
 wire \inv_in[544] ;
 wire \inv_in[545] ;
 wire \inv_in[546] ;
 wire \inv_in[547] ;
 wire \inv_in[548] ;
 wire \inv_in[549] ;
 wire \inv_in[54] ;
 wire \inv_in[550] ;
 wire \inv_in[551] ;
 wire \inv_in[552] ;
 wire \inv_in[553] ;
 wire \inv_in[554] ;
 wire \inv_in[555] ;
 wire \inv_in[556] ;
 wire \inv_in[557] ;
 wire \inv_in[558] ;
 wire \inv_in[559] ;
 wire \inv_in[55] ;
 wire \inv_in[560] ;
 wire \inv_in[561] ;
 wire \inv_in[562] ;
 wire \inv_in[563] ;
 wire \inv_in[564] ;
 wire \inv_in[565] ;
 wire \inv_in[566] ;
 wire \inv_in[567] ;
 wire \inv_in[568] ;
 wire \inv_in[569] ;
 wire \inv_in[56] ;
 wire \inv_in[570] ;
 wire \inv_in[571] ;
 wire \inv_in[572] ;
 wire \inv_in[573] ;
 wire \inv_in[574] ;
 wire \inv_in[575] ;
 wire \inv_in[576] ;
 wire \inv_in[577] ;
 wire \inv_in[578] ;
 wire \inv_in[579] ;
 wire \inv_in[57] ;
 wire \inv_in[580] ;
 wire \inv_in[581] ;
 wire \inv_in[582] ;
 wire \inv_in[583] ;
 wire \inv_in[584] ;
 wire \inv_in[585] ;
 wire \inv_in[586] ;
 wire \inv_in[587] ;
 wire \inv_in[588] ;
 wire \inv_in[589] ;
 wire \inv_in[58] ;
 wire \inv_in[590] ;
 wire \inv_in[591] ;
 wire \inv_in[592] ;
 wire \inv_in[593] ;
 wire \inv_in[594] ;
 wire \inv_in[595] ;
 wire \inv_in[596] ;
 wire \inv_in[597] ;
 wire \inv_in[598] ;
 wire \inv_in[599] ;
 wire \inv_in[59] ;
 wire \inv_in[5] ;
 wire \inv_in[600] ;
 wire \inv_in[601] ;
 wire \inv_in[602] ;
 wire \inv_in[603] ;
 wire \inv_in[604] ;
 wire \inv_in[605] ;
 wire \inv_in[606] ;
 wire \inv_in[607] ;
 wire \inv_in[608] ;
 wire \inv_in[609] ;
 wire \inv_in[60] ;
 wire \inv_in[610] ;
 wire \inv_in[611] ;
 wire \inv_in[612] ;
 wire \inv_in[613] ;
 wire \inv_in[614] ;
 wire \inv_in[615] ;
 wire \inv_in[616] ;
 wire \inv_in[617] ;
 wire \inv_in[618] ;
 wire \inv_in[619] ;
 wire \inv_in[61] ;
 wire \inv_in[620] ;
 wire \inv_in[621] ;
 wire \inv_in[622] ;
 wire \inv_in[623] ;
 wire \inv_in[624] ;
 wire \inv_in[625] ;
 wire \inv_in[626] ;
 wire \inv_in[627] ;
 wire \inv_in[628] ;
 wire \inv_in[629] ;
 wire \inv_in[62] ;
 wire \inv_in[630] ;
 wire \inv_in[631] ;
 wire \inv_in[632] ;
 wire \inv_in[633] ;
 wire \inv_in[634] ;
 wire \inv_in[635] ;
 wire \inv_in[636] ;
 wire \inv_in[637] ;
 wire \inv_in[638] ;
 wire \inv_in[639] ;
 wire \inv_in[63] ;
 wire \inv_in[640] ;
 wire \inv_in[641] ;
 wire \inv_in[642] ;
 wire \inv_in[643] ;
 wire \inv_in[644] ;
 wire \inv_in[645] ;
 wire \inv_in[646] ;
 wire \inv_in[647] ;
 wire \inv_in[648] ;
 wire \inv_in[649] ;
 wire \inv_in[64] ;
 wire \inv_in[650] ;
 wire \inv_in[651] ;
 wire \inv_in[652] ;
 wire \inv_in[653] ;
 wire \inv_in[654] ;
 wire \inv_in[655] ;
 wire \inv_in[656] ;
 wire \inv_in[657] ;
 wire \inv_in[658] ;
 wire \inv_in[659] ;
 wire \inv_in[65] ;
 wire \inv_in[660] ;
 wire \inv_in[661] ;
 wire \inv_in[662] ;
 wire \inv_in[663] ;
 wire \inv_in[664] ;
 wire \inv_in[665] ;
 wire \inv_in[666] ;
 wire \inv_in[667] ;
 wire \inv_in[668] ;
 wire \inv_in[669] ;
 wire \inv_in[66] ;
 wire \inv_in[670] ;
 wire \inv_in[671] ;
 wire \inv_in[672] ;
 wire \inv_in[673] ;
 wire \inv_in[674] ;
 wire \inv_in[675] ;
 wire \inv_in[676] ;
 wire \inv_in[677] ;
 wire \inv_in[678] ;
 wire \inv_in[679] ;
 wire \inv_in[67] ;
 wire \inv_in[680] ;
 wire \inv_in[681] ;
 wire \inv_in[682] ;
 wire \inv_in[683] ;
 wire \inv_in[684] ;
 wire \inv_in[685] ;
 wire \inv_in[686] ;
 wire \inv_in[687] ;
 wire \inv_in[688] ;
 wire \inv_in[689] ;
 wire \inv_in[68] ;
 wire \inv_in[690] ;
 wire \inv_in[691] ;
 wire \inv_in[692] ;
 wire \inv_in[693] ;
 wire \inv_in[694] ;
 wire \inv_in[695] ;
 wire \inv_in[696] ;
 wire \inv_in[697] ;
 wire \inv_in[698] ;
 wire \inv_in[699] ;
 wire \inv_in[69] ;
 wire \inv_in[6] ;
 wire \inv_in[700] ;
 wire \inv_in[701] ;
 wire \inv_in[702] ;
 wire \inv_in[703] ;
 wire \inv_in[704] ;
 wire \inv_in[705] ;
 wire \inv_in[706] ;
 wire \inv_in[707] ;
 wire \inv_in[708] ;
 wire \inv_in[709] ;
 wire \inv_in[70] ;
 wire \inv_in[710] ;
 wire \inv_in[711] ;
 wire \inv_in[712] ;
 wire \inv_in[713] ;
 wire \inv_in[714] ;
 wire \inv_in[715] ;
 wire \inv_in[716] ;
 wire \inv_in[717] ;
 wire \inv_in[718] ;
 wire \inv_in[719] ;
 wire \inv_in[71] ;
 wire \inv_in[720] ;
 wire \inv_in[721] ;
 wire \inv_in[722] ;
 wire \inv_in[723] ;
 wire \inv_in[724] ;
 wire \inv_in[725] ;
 wire \inv_in[726] ;
 wire \inv_in[727] ;
 wire \inv_in[728] ;
 wire \inv_in[729] ;
 wire \inv_in[72] ;
 wire \inv_in[730] ;
 wire \inv_in[731] ;
 wire \inv_in[732] ;
 wire \inv_in[733] ;
 wire \inv_in[734] ;
 wire \inv_in[735] ;
 wire \inv_in[736] ;
 wire \inv_in[737] ;
 wire \inv_in[738] ;
 wire \inv_in[739] ;
 wire \inv_in[73] ;
 wire \inv_in[740] ;
 wire \inv_in[741] ;
 wire \inv_in[742] ;
 wire \inv_in[743] ;
 wire \inv_in[744] ;
 wire \inv_in[745] ;
 wire \inv_in[746] ;
 wire \inv_in[747] ;
 wire \inv_in[748] ;
 wire \inv_in[749] ;
 wire \inv_in[74] ;
 wire \inv_in[750] ;
 wire \inv_in[751] ;
 wire \inv_in[752] ;
 wire \inv_in[753] ;
 wire \inv_in[754] ;
 wire \inv_in[755] ;
 wire \inv_in[756] ;
 wire \inv_in[757] ;
 wire \inv_in[758] ;
 wire \inv_in[759] ;
 wire \inv_in[75] ;
 wire \inv_in[760] ;
 wire \inv_in[761] ;
 wire \inv_in[762] ;
 wire \inv_in[763] ;
 wire \inv_in[764] ;
 wire \inv_in[765] ;
 wire \inv_in[766] ;
 wire \inv_in[767] ;
 wire \inv_in[768] ;
 wire \inv_in[769] ;
 wire \inv_in[76] ;
 wire \inv_in[770] ;
 wire \inv_in[771] ;
 wire \inv_in[772] ;
 wire \inv_in[773] ;
 wire \inv_in[774] ;
 wire \inv_in[775] ;
 wire \inv_in[776] ;
 wire \inv_in[777] ;
 wire \inv_in[778] ;
 wire \inv_in[779] ;
 wire \inv_in[77] ;
 wire \inv_in[780] ;
 wire \inv_in[781] ;
 wire \inv_in[782] ;
 wire \inv_in[783] ;
 wire \inv_in[784] ;
 wire \inv_in[785] ;
 wire \inv_in[786] ;
 wire \inv_in[787] ;
 wire \inv_in[788] ;
 wire \inv_in[789] ;
 wire \inv_in[78] ;
 wire \inv_in[790] ;
 wire \inv_in[791] ;
 wire \inv_in[792] ;
 wire \inv_in[793] ;
 wire \inv_in[794] ;
 wire \inv_in[795] ;
 wire \inv_in[796] ;
 wire \inv_in[797] ;
 wire \inv_in[798] ;
 wire \inv_in[799] ;
 wire \inv_in[79] ;
 wire \inv_in[7] ;
 wire \inv_in[800] ;
 wire \inv_in[801] ;
 wire \inv_in[802] ;
 wire \inv_in[803] ;
 wire \inv_in[804] ;
 wire \inv_in[805] ;
 wire \inv_in[806] ;
 wire \inv_in[807] ;
 wire \inv_in[808] ;
 wire \inv_in[809] ;
 wire \inv_in[80] ;
 wire \inv_in[810] ;
 wire \inv_in[811] ;
 wire \inv_in[812] ;
 wire \inv_in[813] ;
 wire \inv_in[814] ;
 wire \inv_in[815] ;
 wire \inv_in[816] ;
 wire \inv_in[817] ;
 wire \inv_in[818] ;
 wire \inv_in[819] ;
 wire \inv_in[81] ;
 wire \inv_in[820] ;
 wire \inv_in[821] ;
 wire \inv_in[822] ;
 wire \inv_in[823] ;
 wire \inv_in[824] ;
 wire \inv_in[825] ;
 wire \inv_in[826] ;
 wire \inv_in[827] ;
 wire \inv_in[828] ;
 wire \inv_in[829] ;
 wire \inv_in[82] ;
 wire \inv_in[830] ;
 wire \inv_in[831] ;
 wire \inv_in[832] ;
 wire \inv_in[833] ;
 wire \inv_in[834] ;
 wire \inv_in[835] ;
 wire \inv_in[836] ;
 wire \inv_in[837] ;
 wire \inv_in[838] ;
 wire \inv_in[839] ;
 wire \inv_in[83] ;
 wire \inv_in[840] ;
 wire \inv_in[841] ;
 wire \inv_in[842] ;
 wire \inv_in[843] ;
 wire \inv_in[844] ;
 wire \inv_in[845] ;
 wire \inv_in[846] ;
 wire \inv_in[847] ;
 wire \inv_in[848] ;
 wire \inv_in[849] ;
 wire \inv_in[84] ;
 wire \inv_in[850] ;
 wire \inv_in[851] ;
 wire \inv_in[852] ;
 wire \inv_in[853] ;
 wire \inv_in[854] ;
 wire \inv_in[855] ;
 wire \inv_in[856] ;
 wire \inv_in[857] ;
 wire \inv_in[858] ;
 wire \inv_in[859] ;
 wire \inv_in[85] ;
 wire \inv_in[860] ;
 wire \inv_in[861] ;
 wire \inv_in[862] ;
 wire \inv_in[863] ;
 wire \inv_in[864] ;
 wire \inv_in[865] ;
 wire \inv_in[866] ;
 wire \inv_in[867] ;
 wire \inv_in[868] ;
 wire \inv_in[869] ;
 wire \inv_in[86] ;
 wire \inv_in[870] ;
 wire \inv_in[871] ;
 wire \inv_in[872] ;
 wire \inv_in[873] ;
 wire \inv_in[874] ;
 wire \inv_in[875] ;
 wire \inv_in[876] ;
 wire \inv_in[877] ;
 wire \inv_in[878] ;
 wire \inv_in[879] ;
 wire \inv_in[87] ;
 wire \inv_in[880] ;
 wire \inv_in[881] ;
 wire \inv_in[882] ;
 wire \inv_in[883] ;
 wire \inv_in[884] ;
 wire \inv_in[885] ;
 wire \inv_in[886] ;
 wire \inv_in[887] ;
 wire \inv_in[888] ;
 wire \inv_in[889] ;
 wire \inv_in[88] ;
 wire \inv_in[890] ;
 wire \inv_in[891] ;
 wire \inv_in[892] ;
 wire \inv_in[893] ;
 wire \inv_in[894] ;
 wire \inv_in[895] ;
 wire \inv_in[896] ;
 wire \inv_in[897] ;
 wire \inv_in[898] ;
 wire \inv_in[899] ;
 wire \inv_in[89] ;
 wire \inv_in[8] ;
 wire \inv_in[900] ;
 wire \inv_in[901] ;
 wire \inv_in[902] ;
 wire \inv_in[903] ;
 wire \inv_in[904] ;
 wire \inv_in[905] ;
 wire \inv_in[906] ;
 wire \inv_in[907] ;
 wire \inv_in[908] ;
 wire \inv_in[909] ;
 wire \inv_in[90] ;
 wire \inv_in[910] ;
 wire \inv_in[911] ;
 wire \inv_in[912] ;
 wire \inv_in[913] ;
 wire \inv_in[914] ;
 wire \inv_in[915] ;
 wire \inv_in[916] ;
 wire \inv_in[917] ;
 wire \inv_in[918] ;
 wire \inv_in[919] ;
 wire \inv_in[91] ;
 wire \inv_in[920] ;
 wire \inv_in[921] ;
 wire \inv_in[922] ;
 wire \inv_in[923] ;
 wire \inv_in[924] ;
 wire \inv_in[925] ;
 wire \inv_in[926] ;
 wire \inv_in[927] ;
 wire \inv_in[928] ;
 wire \inv_in[929] ;
 wire \inv_in[92] ;
 wire \inv_in[930] ;
 wire \inv_in[931] ;
 wire \inv_in[932] ;
 wire \inv_in[933] ;
 wire \inv_in[934] ;
 wire \inv_in[935] ;
 wire \inv_in[936] ;
 wire \inv_in[937] ;
 wire \inv_in[938] ;
 wire \inv_in[939] ;
 wire \inv_in[93] ;
 wire \inv_in[940] ;
 wire \inv_in[941] ;
 wire \inv_in[942] ;
 wire \inv_in[943] ;
 wire \inv_in[944] ;
 wire \inv_in[945] ;
 wire \inv_in[946] ;
 wire \inv_in[947] ;
 wire \inv_in[948] ;
 wire \inv_in[949] ;
 wire \inv_in[94] ;
 wire \inv_in[950] ;
 wire \inv_in[951] ;
 wire \inv_in[952] ;
 wire \inv_in[953] ;
 wire \inv_in[954] ;
 wire \inv_in[955] ;
 wire \inv_in[956] ;
 wire \inv_in[957] ;
 wire \inv_in[958] ;
 wire \inv_in[959] ;
 wire \inv_in[95] ;
 wire \inv_in[960] ;
 wire \inv_in[961] ;
 wire \inv_in[962] ;
 wire \inv_in[963] ;
 wire \inv_in[964] ;
 wire \inv_in[965] ;
 wire \inv_in[966] ;
 wire \inv_in[967] ;
 wire \inv_in[968] ;
 wire \inv_in[969] ;
 wire \inv_in[96] ;
 wire \inv_in[970] ;
 wire \inv_in[971] ;
 wire \inv_in[972] ;
 wire \inv_in[973] ;
 wire \inv_in[974] ;
 wire \inv_in[975] ;
 wire \inv_in[976] ;
 wire \inv_in[977] ;
 wire \inv_in[978] ;
 wire \inv_in[979] ;
 wire \inv_in[97] ;
 wire \inv_in[980] ;
 wire \inv_in[981] ;
 wire \inv_in[982] ;
 wire \inv_in[983] ;
 wire \inv_in[984] ;
 wire \inv_in[985] ;
 wire \inv_in[986] ;
 wire \inv_in[987] ;
 wire \inv_in[988] ;
 wire \inv_in[989] ;
 wire \inv_in[98] ;
 wire \inv_in[990] ;
 wire \inv_in[991] ;
 wire \inv_in[992] ;
 wire \inv_in[993] ;
 wire \inv_in[994] ;
 wire \inv_in[995] ;
 wire \inv_in[996] ;
 wire \inv_in[997] ;
 wire \inv_in[998] ;
 wire \inv_in[999] ;
 wire \inv_in[99] ;
 wire \inv_in[9] ;
 wire net10;
 wire net11;
 wire net12;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net4;
 wire net5;
 wire net1;
 wire net2;
 wire net3;

 sky130_fd_sc_hd__mux2_1 _00_ (.A0(net1),
    .A1(uio_out[5]),
    .S(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\inv_in[0] ));
 sky130_fd_sc_hd__conb_1 tt_um_urish_giant_ringosc_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net6));
 sky130_fd_sc_hd__conb_1 tt_um_urish_giant_ringosc_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net7));
 sky130_fd_sc_hd__conb_1 tt_um_urish_giant_ringosc_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net8));
 sky130_fd_sc_hd__conb_1 tt_um_urish_giant_ringosc_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net9));
 sky130_fd_sc_hd__conb_1 tt_um_urish_giant_ringosc_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net10));
 sky130_fd_sc_hd__conb_1 tt_um_urish_giant_ringosc_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net11));
 sky130_fd_sc_hd__conb_1 tt_um_urish_giant_ringosc_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net12));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 tt_um_urish_giant_ringosc_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net4));
 sky130_fd_sc_hd__conb_1 tt_um_urish_giant_ringosc_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net5));
 sky130_fd_sc_hd__buf_2 _11_ (.A(\inv_in[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[0]));
 sky130_fd_sc_hd__buf_2 _12_ (.A(\inv_in[501] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[1]));
 sky130_fd_sc_hd__buf_2 _13_ (.A(\inv_in[1001] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[2]));
 sky130_fd_sc_hd__buf_2 _14_ (.A(\inv_in[2001] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[3]));
 sky130_fd_sc_hd__buf_2 _15_ (.A(\inv_in[3001] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__buf_2 _16_ (.A(\inv_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _17_ (.A(\inv_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__buf_2 _18_ (.A(\inv_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__buf_2 _19_ (.A(\inv_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__buf_2 _20_ (.A(\inv_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__buf_2 _21_ (.A(\inv_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__buf_2 _22_ (.A(\inv_in[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__buf_2 _23_ (.A(\inv_in[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__inv_2 \inv[0]/_0_  (.A(\inv_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1] ));
 sky130_fd_sc_hd__inv_2 \inv[1000]/_0_  (.A(\inv_in[1000] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1001] ));
 sky130_fd_sc_hd__inv_2 \inv[1001]/_0_  (.A(\inv_in[1001] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1002] ));
 sky130_fd_sc_hd__inv_2 \inv[1002]/_0_  (.A(\inv_in[1002] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1003] ));
 sky130_fd_sc_hd__inv_2 \inv[1003]/_0_  (.A(\inv_in[1003] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1004] ));
 sky130_fd_sc_hd__inv_2 \inv[1004]/_0_  (.A(\inv_in[1004] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1005] ));
 sky130_fd_sc_hd__inv_2 \inv[1005]/_0_  (.A(\inv_in[1005] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1006] ));
 sky130_fd_sc_hd__inv_2 \inv[1006]/_0_  (.A(\inv_in[1006] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1007] ));
 sky130_fd_sc_hd__inv_2 \inv[1007]/_0_  (.A(\inv_in[1007] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1008] ));
 sky130_fd_sc_hd__inv_2 \inv[1008]/_0_  (.A(\inv_in[1008] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1009] ));
 sky130_fd_sc_hd__inv_2 \inv[1009]/_0_  (.A(\inv_in[1009] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1010] ));
 sky130_fd_sc_hd__inv_2 \inv[100]/_0_  (.A(\inv_in[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[101] ));
 sky130_fd_sc_hd__inv_2 \inv[1010]/_0_  (.A(\inv_in[1010] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1011] ));
 sky130_fd_sc_hd__inv_2 \inv[1011]/_0_  (.A(\inv_in[1011] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1012] ));
 sky130_fd_sc_hd__inv_2 \inv[1012]/_0_  (.A(\inv_in[1012] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1013] ));
 sky130_fd_sc_hd__inv_2 \inv[1013]/_0_  (.A(\inv_in[1013] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1014] ));
 sky130_fd_sc_hd__inv_2 \inv[1014]/_0_  (.A(\inv_in[1014] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1015] ));
 sky130_fd_sc_hd__inv_2 \inv[1015]/_0_  (.A(\inv_in[1015] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1016] ));
 sky130_fd_sc_hd__inv_2 \inv[1016]/_0_  (.A(\inv_in[1016] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1017] ));
 sky130_fd_sc_hd__inv_2 \inv[1017]/_0_  (.A(\inv_in[1017] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1018] ));
 sky130_fd_sc_hd__inv_2 \inv[1018]/_0_  (.A(\inv_in[1018] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1019] ));
 sky130_fd_sc_hd__inv_2 \inv[1019]/_0_  (.A(\inv_in[1019] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1020] ));
 sky130_fd_sc_hd__inv_2 \inv[101]/_0_  (.A(\inv_in[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[102] ));
 sky130_fd_sc_hd__inv_2 \inv[1020]/_0_  (.A(\inv_in[1020] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1021] ));
 sky130_fd_sc_hd__inv_2 \inv[1021]/_0_  (.A(\inv_in[1021] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1022] ));
 sky130_fd_sc_hd__inv_2 \inv[1022]/_0_  (.A(\inv_in[1022] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1023] ));
 sky130_fd_sc_hd__inv_2 \inv[1023]/_0_  (.A(\inv_in[1023] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1024] ));
 sky130_fd_sc_hd__inv_2 \inv[1024]/_0_  (.A(\inv_in[1024] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1025] ));
 sky130_fd_sc_hd__inv_2 \inv[1025]/_0_  (.A(\inv_in[1025] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1026] ));
 sky130_fd_sc_hd__inv_2 \inv[1026]/_0_  (.A(\inv_in[1026] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1027] ));
 sky130_fd_sc_hd__inv_2 \inv[1027]/_0_  (.A(\inv_in[1027] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1028] ));
 sky130_fd_sc_hd__inv_2 \inv[1028]/_0_  (.A(\inv_in[1028] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1029] ));
 sky130_fd_sc_hd__inv_2 \inv[1029]/_0_  (.A(\inv_in[1029] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1030] ));
 sky130_fd_sc_hd__inv_2 \inv[102]/_0_  (.A(\inv_in[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[103] ));
 sky130_fd_sc_hd__inv_2 \inv[1030]/_0_  (.A(\inv_in[1030] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1031] ));
 sky130_fd_sc_hd__inv_2 \inv[1031]/_0_  (.A(\inv_in[1031] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1032] ));
 sky130_fd_sc_hd__inv_2 \inv[1032]/_0_  (.A(\inv_in[1032] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1033] ));
 sky130_fd_sc_hd__inv_2 \inv[1033]/_0_  (.A(\inv_in[1033] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1034] ));
 sky130_fd_sc_hd__inv_2 \inv[1034]/_0_  (.A(\inv_in[1034] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1035] ));
 sky130_fd_sc_hd__inv_2 \inv[1035]/_0_  (.A(\inv_in[1035] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1036] ));
 sky130_fd_sc_hd__inv_2 \inv[1036]/_0_  (.A(\inv_in[1036] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1037] ));
 sky130_fd_sc_hd__inv_2 \inv[1037]/_0_  (.A(\inv_in[1037] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1038] ));
 sky130_fd_sc_hd__inv_2 \inv[1038]/_0_  (.A(\inv_in[1038] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1039] ));
 sky130_fd_sc_hd__inv_2 \inv[1039]/_0_  (.A(\inv_in[1039] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1040] ));
 sky130_fd_sc_hd__inv_2 \inv[103]/_0_  (.A(\inv_in[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[104] ));
 sky130_fd_sc_hd__inv_2 \inv[1040]/_0_  (.A(\inv_in[1040] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1041] ));
 sky130_fd_sc_hd__inv_2 \inv[1041]/_0_  (.A(\inv_in[1041] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1042] ));
 sky130_fd_sc_hd__inv_2 \inv[1042]/_0_  (.A(\inv_in[1042] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1043] ));
 sky130_fd_sc_hd__inv_2 \inv[1043]/_0_  (.A(\inv_in[1043] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1044] ));
 sky130_fd_sc_hd__inv_2 \inv[1044]/_0_  (.A(\inv_in[1044] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1045] ));
 sky130_fd_sc_hd__inv_2 \inv[1045]/_0_  (.A(\inv_in[1045] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1046] ));
 sky130_fd_sc_hd__inv_2 \inv[1046]/_0_  (.A(\inv_in[1046] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1047] ));
 sky130_fd_sc_hd__inv_2 \inv[1047]/_0_  (.A(\inv_in[1047] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1048] ));
 sky130_fd_sc_hd__inv_2 \inv[1048]/_0_  (.A(\inv_in[1048] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1049] ));
 sky130_fd_sc_hd__inv_2 \inv[1049]/_0_  (.A(\inv_in[1049] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1050] ));
 sky130_fd_sc_hd__inv_2 \inv[104]/_0_  (.A(\inv_in[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[105] ));
 sky130_fd_sc_hd__inv_2 \inv[1050]/_0_  (.A(\inv_in[1050] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1051] ));
 sky130_fd_sc_hd__inv_2 \inv[1051]/_0_  (.A(\inv_in[1051] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1052] ));
 sky130_fd_sc_hd__inv_2 \inv[1052]/_0_  (.A(\inv_in[1052] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1053] ));
 sky130_fd_sc_hd__inv_2 \inv[1053]/_0_  (.A(\inv_in[1053] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1054] ));
 sky130_fd_sc_hd__inv_2 \inv[1054]/_0_  (.A(\inv_in[1054] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1055] ));
 sky130_fd_sc_hd__inv_2 \inv[1055]/_0_  (.A(\inv_in[1055] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1056] ));
 sky130_fd_sc_hd__inv_2 \inv[1056]/_0_  (.A(\inv_in[1056] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1057] ));
 sky130_fd_sc_hd__inv_2 \inv[1057]/_0_  (.A(\inv_in[1057] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1058] ));
 sky130_fd_sc_hd__inv_2 \inv[1058]/_0_  (.A(\inv_in[1058] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1059] ));
 sky130_fd_sc_hd__inv_2 \inv[1059]/_0_  (.A(\inv_in[1059] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1060] ));
 sky130_fd_sc_hd__inv_2 \inv[105]/_0_  (.A(\inv_in[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[106] ));
 sky130_fd_sc_hd__inv_2 \inv[1060]/_0_  (.A(\inv_in[1060] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1061] ));
 sky130_fd_sc_hd__inv_2 \inv[1061]/_0_  (.A(\inv_in[1061] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1062] ));
 sky130_fd_sc_hd__inv_2 \inv[1062]/_0_  (.A(\inv_in[1062] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1063] ));
 sky130_fd_sc_hd__inv_2 \inv[1063]/_0_  (.A(\inv_in[1063] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1064] ));
 sky130_fd_sc_hd__inv_2 \inv[1064]/_0_  (.A(\inv_in[1064] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1065] ));
 sky130_fd_sc_hd__inv_2 \inv[1065]/_0_  (.A(\inv_in[1065] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1066] ));
 sky130_fd_sc_hd__inv_2 \inv[1066]/_0_  (.A(\inv_in[1066] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1067] ));
 sky130_fd_sc_hd__inv_2 \inv[1067]/_0_  (.A(\inv_in[1067] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1068] ));
 sky130_fd_sc_hd__inv_2 \inv[1068]/_0_  (.A(\inv_in[1068] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1069] ));
 sky130_fd_sc_hd__inv_2 \inv[1069]/_0_  (.A(\inv_in[1069] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1070] ));
 sky130_fd_sc_hd__inv_2 \inv[106]/_0_  (.A(\inv_in[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[107] ));
 sky130_fd_sc_hd__inv_2 \inv[1070]/_0_  (.A(\inv_in[1070] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1071] ));
 sky130_fd_sc_hd__inv_2 \inv[1071]/_0_  (.A(\inv_in[1071] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1072] ));
 sky130_fd_sc_hd__inv_2 \inv[1072]/_0_  (.A(\inv_in[1072] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1073] ));
 sky130_fd_sc_hd__inv_2 \inv[1073]/_0_  (.A(\inv_in[1073] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1074] ));
 sky130_fd_sc_hd__inv_2 \inv[1074]/_0_  (.A(\inv_in[1074] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1075] ));
 sky130_fd_sc_hd__inv_2 \inv[1075]/_0_  (.A(\inv_in[1075] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1076] ));
 sky130_fd_sc_hd__inv_2 \inv[1076]/_0_  (.A(\inv_in[1076] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1077] ));
 sky130_fd_sc_hd__inv_2 \inv[1077]/_0_  (.A(\inv_in[1077] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1078] ));
 sky130_fd_sc_hd__inv_2 \inv[1078]/_0_  (.A(\inv_in[1078] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1079] ));
 sky130_fd_sc_hd__inv_2 \inv[1079]/_0_  (.A(\inv_in[1079] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1080] ));
 sky130_fd_sc_hd__inv_2 \inv[107]/_0_  (.A(\inv_in[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[108] ));
 sky130_fd_sc_hd__inv_2 \inv[1080]/_0_  (.A(\inv_in[1080] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1081] ));
 sky130_fd_sc_hd__inv_2 \inv[1081]/_0_  (.A(\inv_in[1081] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1082] ));
 sky130_fd_sc_hd__inv_2 \inv[1082]/_0_  (.A(\inv_in[1082] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1083] ));
 sky130_fd_sc_hd__inv_2 \inv[1083]/_0_  (.A(\inv_in[1083] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1084] ));
 sky130_fd_sc_hd__inv_2 \inv[1084]/_0_  (.A(\inv_in[1084] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1085] ));
 sky130_fd_sc_hd__inv_2 \inv[1085]/_0_  (.A(\inv_in[1085] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1086] ));
 sky130_fd_sc_hd__inv_2 \inv[1086]/_0_  (.A(\inv_in[1086] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1087] ));
 sky130_fd_sc_hd__inv_2 \inv[1087]/_0_  (.A(\inv_in[1087] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1088] ));
 sky130_fd_sc_hd__inv_2 \inv[1088]/_0_  (.A(\inv_in[1088] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1089] ));
 sky130_fd_sc_hd__inv_2 \inv[1089]/_0_  (.A(\inv_in[1089] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1090] ));
 sky130_fd_sc_hd__inv_2 \inv[108]/_0_  (.A(\inv_in[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[109] ));
 sky130_fd_sc_hd__inv_2 \inv[1090]/_0_  (.A(\inv_in[1090] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1091] ));
 sky130_fd_sc_hd__inv_2 \inv[1091]/_0_  (.A(\inv_in[1091] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1092] ));
 sky130_fd_sc_hd__inv_2 \inv[1092]/_0_  (.A(\inv_in[1092] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1093] ));
 sky130_fd_sc_hd__inv_2 \inv[1093]/_0_  (.A(\inv_in[1093] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1094] ));
 sky130_fd_sc_hd__inv_2 \inv[1094]/_0_  (.A(\inv_in[1094] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1095] ));
 sky130_fd_sc_hd__inv_2 \inv[1095]/_0_  (.A(\inv_in[1095] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1096] ));
 sky130_fd_sc_hd__inv_2 \inv[1096]/_0_  (.A(\inv_in[1096] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1097] ));
 sky130_fd_sc_hd__inv_2 \inv[1097]/_0_  (.A(\inv_in[1097] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1098] ));
 sky130_fd_sc_hd__inv_2 \inv[1098]/_0_  (.A(\inv_in[1098] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1099] ));
 sky130_fd_sc_hd__inv_2 \inv[1099]/_0_  (.A(\inv_in[1099] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1100] ));
 sky130_fd_sc_hd__inv_2 \inv[109]/_0_  (.A(\inv_in[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[110] ));
 sky130_fd_sc_hd__inv_2 \inv[10]/_0_  (.A(\inv_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[11] ));
 sky130_fd_sc_hd__inv_2 \inv[1100]/_0_  (.A(\inv_in[1100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1101] ));
 sky130_fd_sc_hd__inv_2 \inv[1101]/_0_  (.A(\inv_in[1101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1102] ));
 sky130_fd_sc_hd__inv_2 \inv[1102]/_0_  (.A(\inv_in[1102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1103] ));
 sky130_fd_sc_hd__inv_2 \inv[1103]/_0_  (.A(\inv_in[1103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1104] ));
 sky130_fd_sc_hd__inv_2 \inv[1104]/_0_  (.A(\inv_in[1104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1105] ));
 sky130_fd_sc_hd__inv_2 \inv[1105]/_0_  (.A(\inv_in[1105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1106] ));
 sky130_fd_sc_hd__inv_2 \inv[1106]/_0_  (.A(\inv_in[1106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1107] ));
 sky130_fd_sc_hd__inv_2 \inv[1107]/_0_  (.A(\inv_in[1107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1108] ));
 sky130_fd_sc_hd__inv_2 \inv[1108]/_0_  (.A(\inv_in[1108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1109] ));
 sky130_fd_sc_hd__inv_2 \inv[1109]/_0_  (.A(\inv_in[1109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1110] ));
 sky130_fd_sc_hd__inv_2 \inv[110]/_0_  (.A(\inv_in[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[111] ));
 sky130_fd_sc_hd__inv_2 \inv[1110]/_0_  (.A(\inv_in[1110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1111] ));
 sky130_fd_sc_hd__inv_2 \inv[1111]/_0_  (.A(\inv_in[1111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1112] ));
 sky130_fd_sc_hd__inv_2 \inv[1112]/_0_  (.A(\inv_in[1112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1113] ));
 sky130_fd_sc_hd__inv_2 \inv[1113]/_0_  (.A(\inv_in[1113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1114] ));
 sky130_fd_sc_hd__inv_2 \inv[1114]/_0_  (.A(\inv_in[1114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1115] ));
 sky130_fd_sc_hd__inv_2 \inv[1115]/_0_  (.A(\inv_in[1115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1116] ));
 sky130_fd_sc_hd__inv_2 \inv[1116]/_0_  (.A(\inv_in[1116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1117] ));
 sky130_fd_sc_hd__inv_2 \inv[1117]/_0_  (.A(\inv_in[1117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1118] ));
 sky130_fd_sc_hd__inv_2 \inv[1118]/_0_  (.A(\inv_in[1118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1119] ));
 sky130_fd_sc_hd__inv_2 \inv[1119]/_0_  (.A(\inv_in[1119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1120] ));
 sky130_fd_sc_hd__inv_2 \inv[111]/_0_  (.A(\inv_in[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[112] ));
 sky130_fd_sc_hd__inv_2 \inv[1120]/_0_  (.A(\inv_in[1120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1121] ));
 sky130_fd_sc_hd__inv_2 \inv[1121]/_0_  (.A(\inv_in[1121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1122] ));
 sky130_fd_sc_hd__inv_2 \inv[1122]/_0_  (.A(\inv_in[1122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1123] ));
 sky130_fd_sc_hd__inv_2 \inv[1123]/_0_  (.A(\inv_in[1123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1124] ));
 sky130_fd_sc_hd__inv_2 \inv[1124]/_0_  (.A(\inv_in[1124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1125] ));
 sky130_fd_sc_hd__inv_2 \inv[1125]/_0_  (.A(\inv_in[1125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1126] ));
 sky130_fd_sc_hd__inv_2 \inv[1126]/_0_  (.A(\inv_in[1126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1127] ));
 sky130_fd_sc_hd__inv_2 \inv[1127]/_0_  (.A(\inv_in[1127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1128] ));
 sky130_fd_sc_hd__inv_2 \inv[1128]/_0_  (.A(\inv_in[1128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1129] ));
 sky130_fd_sc_hd__inv_2 \inv[1129]/_0_  (.A(\inv_in[1129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1130] ));
 sky130_fd_sc_hd__inv_2 \inv[112]/_0_  (.A(\inv_in[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[113] ));
 sky130_fd_sc_hd__inv_2 \inv[1130]/_0_  (.A(\inv_in[1130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1131] ));
 sky130_fd_sc_hd__inv_2 \inv[1131]/_0_  (.A(\inv_in[1131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1132] ));
 sky130_fd_sc_hd__inv_2 \inv[1132]/_0_  (.A(\inv_in[1132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1133] ));
 sky130_fd_sc_hd__inv_2 \inv[1133]/_0_  (.A(\inv_in[1133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1134] ));
 sky130_fd_sc_hd__inv_2 \inv[1134]/_0_  (.A(\inv_in[1134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1135] ));
 sky130_fd_sc_hd__inv_2 \inv[1135]/_0_  (.A(\inv_in[1135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1136] ));
 sky130_fd_sc_hd__inv_2 \inv[1136]/_0_  (.A(\inv_in[1136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1137] ));
 sky130_fd_sc_hd__inv_2 \inv[1137]/_0_  (.A(\inv_in[1137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1138] ));
 sky130_fd_sc_hd__inv_2 \inv[1138]/_0_  (.A(\inv_in[1138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1139] ));
 sky130_fd_sc_hd__inv_2 \inv[1139]/_0_  (.A(\inv_in[1139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1140] ));
 sky130_fd_sc_hd__inv_2 \inv[113]/_0_  (.A(\inv_in[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[114] ));
 sky130_fd_sc_hd__inv_2 \inv[1140]/_0_  (.A(\inv_in[1140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1141] ));
 sky130_fd_sc_hd__inv_2 \inv[1141]/_0_  (.A(\inv_in[1141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1142] ));
 sky130_fd_sc_hd__inv_2 \inv[1142]/_0_  (.A(\inv_in[1142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1143] ));
 sky130_fd_sc_hd__inv_2 \inv[1143]/_0_  (.A(\inv_in[1143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1144] ));
 sky130_fd_sc_hd__inv_2 \inv[1144]/_0_  (.A(\inv_in[1144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1145] ));
 sky130_fd_sc_hd__inv_2 \inv[1145]/_0_  (.A(\inv_in[1145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1146] ));
 sky130_fd_sc_hd__inv_2 \inv[1146]/_0_  (.A(\inv_in[1146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1147] ));
 sky130_fd_sc_hd__inv_2 \inv[1147]/_0_  (.A(\inv_in[1147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1148] ));
 sky130_fd_sc_hd__inv_2 \inv[1148]/_0_  (.A(\inv_in[1148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1149] ));
 sky130_fd_sc_hd__inv_2 \inv[1149]/_0_  (.A(\inv_in[1149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1150] ));
 sky130_fd_sc_hd__inv_2 \inv[114]/_0_  (.A(\inv_in[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[115] ));
 sky130_fd_sc_hd__inv_2 \inv[1150]/_0_  (.A(\inv_in[1150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1151] ));
 sky130_fd_sc_hd__inv_2 \inv[1151]/_0_  (.A(\inv_in[1151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1152] ));
 sky130_fd_sc_hd__inv_2 \inv[1152]/_0_  (.A(\inv_in[1152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1153] ));
 sky130_fd_sc_hd__inv_2 \inv[1153]/_0_  (.A(\inv_in[1153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1154] ));
 sky130_fd_sc_hd__inv_2 \inv[1154]/_0_  (.A(\inv_in[1154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1155] ));
 sky130_fd_sc_hd__inv_2 \inv[1155]/_0_  (.A(\inv_in[1155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1156] ));
 sky130_fd_sc_hd__inv_2 \inv[1156]/_0_  (.A(\inv_in[1156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1157] ));
 sky130_fd_sc_hd__inv_2 \inv[1157]/_0_  (.A(\inv_in[1157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1158] ));
 sky130_fd_sc_hd__inv_2 \inv[1158]/_0_  (.A(\inv_in[1158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1159] ));
 sky130_fd_sc_hd__inv_2 \inv[1159]/_0_  (.A(\inv_in[1159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1160] ));
 sky130_fd_sc_hd__inv_2 \inv[115]/_0_  (.A(\inv_in[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[116] ));
 sky130_fd_sc_hd__inv_2 \inv[1160]/_0_  (.A(\inv_in[1160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1161] ));
 sky130_fd_sc_hd__inv_2 \inv[1161]/_0_  (.A(\inv_in[1161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1162] ));
 sky130_fd_sc_hd__inv_2 \inv[1162]/_0_  (.A(\inv_in[1162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1163] ));
 sky130_fd_sc_hd__inv_2 \inv[1163]/_0_  (.A(\inv_in[1163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1164] ));
 sky130_fd_sc_hd__inv_2 \inv[1164]/_0_  (.A(\inv_in[1164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1165] ));
 sky130_fd_sc_hd__inv_2 \inv[1165]/_0_  (.A(\inv_in[1165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1166] ));
 sky130_fd_sc_hd__inv_2 \inv[1166]/_0_  (.A(\inv_in[1166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1167] ));
 sky130_fd_sc_hd__inv_2 \inv[1167]/_0_  (.A(\inv_in[1167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1168] ));
 sky130_fd_sc_hd__inv_2 \inv[1168]/_0_  (.A(\inv_in[1168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1169] ));
 sky130_fd_sc_hd__inv_2 \inv[1169]/_0_  (.A(\inv_in[1169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1170] ));
 sky130_fd_sc_hd__inv_2 \inv[116]/_0_  (.A(\inv_in[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[117] ));
 sky130_fd_sc_hd__inv_2 \inv[1170]/_0_  (.A(\inv_in[1170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1171] ));
 sky130_fd_sc_hd__inv_2 \inv[1171]/_0_  (.A(\inv_in[1171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1172] ));
 sky130_fd_sc_hd__inv_2 \inv[1172]/_0_  (.A(\inv_in[1172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1173] ));
 sky130_fd_sc_hd__inv_2 \inv[1173]/_0_  (.A(\inv_in[1173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1174] ));
 sky130_fd_sc_hd__inv_2 \inv[1174]/_0_  (.A(\inv_in[1174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1175] ));
 sky130_fd_sc_hd__inv_2 \inv[1175]/_0_  (.A(\inv_in[1175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1176] ));
 sky130_fd_sc_hd__inv_2 \inv[1176]/_0_  (.A(\inv_in[1176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1177] ));
 sky130_fd_sc_hd__inv_2 \inv[1177]/_0_  (.A(\inv_in[1177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1178] ));
 sky130_fd_sc_hd__inv_2 \inv[1178]/_0_  (.A(\inv_in[1178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1179] ));
 sky130_fd_sc_hd__inv_2 \inv[1179]/_0_  (.A(\inv_in[1179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1180] ));
 sky130_fd_sc_hd__inv_2 \inv[117]/_0_  (.A(\inv_in[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[118] ));
 sky130_fd_sc_hd__inv_2 \inv[1180]/_0_  (.A(\inv_in[1180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1181] ));
 sky130_fd_sc_hd__inv_2 \inv[1181]/_0_  (.A(\inv_in[1181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1182] ));
 sky130_fd_sc_hd__inv_2 \inv[1182]/_0_  (.A(\inv_in[1182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1183] ));
 sky130_fd_sc_hd__inv_2 \inv[1183]/_0_  (.A(\inv_in[1183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1184] ));
 sky130_fd_sc_hd__inv_2 \inv[1184]/_0_  (.A(\inv_in[1184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1185] ));
 sky130_fd_sc_hd__inv_2 \inv[1185]/_0_  (.A(\inv_in[1185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1186] ));
 sky130_fd_sc_hd__inv_2 \inv[1186]/_0_  (.A(\inv_in[1186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1187] ));
 sky130_fd_sc_hd__inv_2 \inv[1187]/_0_  (.A(\inv_in[1187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1188] ));
 sky130_fd_sc_hd__inv_2 \inv[1188]/_0_  (.A(\inv_in[1188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1189] ));
 sky130_fd_sc_hd__inv_2 \inv[1189]/_0_  (.A(\inv_in[1189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1190] ));
 sky130_fd_sc_hd__inv_2 \inv[118]/_0_  (.A(\inv_in[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[119] ));
 sky130_fd_sc_hd__inv_2 \inv[1190]/_0_  (.A(\inv_in[1190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1191] ));
 sky130_fd_sc_hd__inv_2 \inv[1191]/_0_  (.A(\inv_in[1191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1192] ));
 sky130_fd_sc_hd__inv_2 \inv[1192]/_0_  (.A(\inv_in[1192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1193] ));
 sky130_fd_sc_hd__inv_2 \inv[1193]/_0_  (.A(\inv_in[1193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1194] ));
 sky130_fd_sc_hd__inv_2 \inv[1194]/_0_  (.A(\inv_in[1194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1195] ));
 sky130_fd_sc_hd__inv_2 \inv[1195]/_0_  (.A(\inv_in[1195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1196] ));
 sky130_fd_sc_hd__inv_2 \inv[1196]/_0_  (.A(\inv_in[1196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1197] ));
 sky130_fd_sc_hd__inv_2 \inv[1197]/_0_  (.A(\inv_in[1197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1198] ));
 sky130_fd_sc_hd__inv_2 \inv[1198]/_0_  (.A(\inv_in[1198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1199] ));
 sky130_fd_sc_hd__inv_2 \inv[1199]/_0_  (.A(\inv_in[1199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1200] ));
 sky130_fd_sc_hd__inv_2 \inv[119]/_0_  (.A(\inv_in[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[120] ));
 sky130_fd_sc_hd__inv_2 \inv[11]/_0_  (.A(\inv_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[12] ));
 sky130_fd_sc_hd__inv_2 \inv[1200]/_0_  (.A(\inv_in[1200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1201] ));
 sky130_fd_sc_hd__inv_2 \inv[1201]/_0_  (.A(\inv_in[1201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1202] ));
 sky130_fd_sc_hd__inv_2 \inv[1202]/_0_  (.A(\inv_in[1202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1203] ));
 sky130_fd_sc_hd__inv_2 \inv[1203]/_0_  (.A(\inv_in[1203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1204] ));
 sky130_fd_sc_hd__inv_2 \inv[1204]/_0_  (.A(\inv_in[1204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1205] ));
 sky130_fd_sc_hd__inv_2 \inv[1205]/_0_  (.A(\inv_in[1205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1206] ));
 sky130_fd_sc_hd__inv_2 \inv[1206]/_0_  (.A(\inv_in[1206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1207] ));
 sky130_fd_sc_hd__inv_2 \inv[1207]/_0_  (.A(\inv_in[1207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1208] ));
 sky130_fd_sc_hd__inv_2 \inv[1208]/_0_  (.A(\inv_in[1208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1209] ));
 sky130_fd_sc_hd__inv_2 \inv[1209]/_0_  (.A(\inv_in[1209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1210] ));
 sky130_fd_sc_hd__inv_2 \inv[120]/_0_  (.A(\inv_in[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[121] ));
 sky130_fd_sc_hd__inv_2 \inv[1210]/_0_  (.A(\inv_in[1210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1211] ));
 sky130_fd_sc_hd__inv_2 \inv[1211]/_0_  (.A(\inv_in[1211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1212] ));
 sky130_fd_sc_hd__inv_2 \inv[1212]/_0_  (.A(\inv_in[1212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1213] ));
 sky130_fd_sc_hd__inv_2 \inv[1213]/_0_  (.A(\inv_in[1213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1214] ));
 sky130_fd_sc_hd__inv_2 \inv[1214]/_0_  (.A(\inv_in[1214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1215] ));
 sky130_fd_sc_hd__inv_2 \inv[1215]/_0_  (.A(\inv_in[1215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1216] ));
 sky130_fd_sc_hd__inv_2 \inv[1216]/_0_  (.A(\inv_in[1216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1217] ));
 sky130_fd_sc_hd__inv_2 \inv[1217]/_0_  (.A(\inv_in[1217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1218] ));
 sky130_fd_sc_hd__inv_2 \inv[1218]/_0_  (.A(\inv_in[1218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1219] ));
 sky130_fd_sc_hd__inv_2 \inv[1219]/_0_  (.A(\inv_in[1219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1220] ));
 sky130_fd_sc_hd__inv_2 \inv[121]/_0_  (.A(\inv_in[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[122] ));
 sky130_fd_sc_hd__inv_2 \inv[1220]/_0_  (.A(\inv_in[1220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1221] ));
 sky130_fd_sc_hd__inv_2 \inv[1221]/_0_  (.A(\inv_in[1221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1222] ));
 sky130_fd_sc_hd__inv_2 \inv[1222]/_0_  (.A(\inv_in[1222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1223] ));
 sky130_fd_sc_hd__inv_2 \inv[1223]/_0_  (.A(\inv_in[1223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1224] ));
 sky130_fd_sc_hd__inv_2 \inv[1224]/_0_  (.A(\inv_in[1224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1225] ));
 sky130_fd_sc_hd__inv_2 \inv[1225]/_0_  (.A(\inv_in[1225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1226] ));
 sky130_fd_sc_hd__inv_2 \inv[1226]/_0_  (.A(\inv_in[1226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1227] ));
 sky130_fd_sc_hd__inv_2 \inv[1227]/_0_  (.A(\inv_in[1227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1228] ));
 sky130_fd_sc_hd__inv_2 \inv[1228]/_0_  (.A(\inv_in[1228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1229] ));
 sky130_fd_sc_hd__inv_2 \inv[1229]/_0_  (.A(\inv_in[1229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1230] ));
 sky130_fd_sc_hd__inv_2 \inv[122]/_0_  (.A(\inv_in[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[123] ));
 sky130_fd_sc_hd__inv_2 \inv[1230]/_0_  (.A(\inv_in[1230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1231] ));
 sky130_fd_sc_hd__inv_2 \inv[1231]/_0_  (.A(\inv_in[1231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1232] ));
 sky130_fd_sc_hd__inv_2 \inv[1232]/_0_  (.A(\inv_in[1232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1233] ));
 sky130_fd_sc_hd__inv_2 \inv[1233]/_0_  (.A(\inv_in[1233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1234] ));
 sky130_fd_sc_hd__inv_2 \inv[1234]/_0_  (.A(\inv_in[1234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1235] ));
 sky130_fd_sc_hd__inv_2 \inv[1235]/_0_  (.A(\inv_in[1235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1236] ));
 sky130_fd_sc_hd__inv_2 \inv[1236]/_0_  (.A(\inv_in[1236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1237] ));
 sky130_fd_sc_hd__inv_2 \inv[1237]/_0_  (.A(\inv_in[1237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1238] ));
 sky130_fd_sc_hd__inv_2 \inv[1238]/_0_  (.A(\inv_in[1238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1239] ));
 sky130_fd_sc_hd__inv_2 \inv[1239]/_0_  (.A(\inv_in[1239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1240] ));
 sky130_fd_sc_hd__inv_2 \inv[123]/_0_  (.A(\inv_in[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[124] ));
 sky130_fd_sc_hd__inv_2 \inv[1240]/_0_  (.A(\inv_in[1240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1241] ));
 sky130_fd_sc_hd__inv_2 \inv[1241]/_0_  (.A(\inv_in[1241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1242] ));
 sky130_fd_sc_hd__inv_2 \inv[1242]/_0_  (.A(\inv_in[1242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1243] ));
 sky130_fd_sc_hd__inv_2 \inv[1243]/_0_  (.A(\inv_in[1243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1244] ));
 sky130_fd_sc_hd__inv_2 \inv[1244]/_0_  (.A(\inv_in[1244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1245] ));
 sky130_fd_sc_hd__inv_2 \inv[1245]/_0_  (.A(\inv_in[1245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1246] ));
 sky130_fd_sc_hd__inv_2 \inv[1246]/_0_  (.A(\inv_in[1246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1247] ));
 sky130_fd_sc_hd__inv_2 \inv[1247]/_0_  (.A(\inv_in[1247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1248] ));
 sky130_fd_sc_hd__inv_2 \inv[1248]/_0_  (.A(\inv_in[1248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1249] ));
 sky130_fd_sc_hd__inv_2 \inv[1249]/_0_  (.A(\inv_in[1249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1250] ));
 sky130_fd_sc_hd__inv_2 \inv[124]/_0_  (.A(\inv_in[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[125] ));
 sky130_fd_sc_hd__inv_2 \inv[1250]/_0_  (.A(\inv_in[1250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1251] ));
 sky130_fd_sc_hd__inv_2 \inv[1251]/_0_  (.A(\inv_in[1251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1252] ));
 sky130_fd_sc_hd__inv_2 \inv[1252]/_0_  (.A(\inv_in[1252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1253] ));
 sky130_fd_sc_hd__inv_2 \inv[1253]/_0_  (.A(\inv_in[1253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1254] ));
 sky130_fd_sc_hd__inv_2 \inv[1254]/_0_  (.A(\inv_in[1254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1255] ));
 sky130_fd_sc_hd__inv_2 \inv[1255]/_0_  (.A(\inv_in[1255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1256] ));
 sky130_fd_sc_hd__inv_2 \inv[1256]/_0_  (.A(\inv_in[1256] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1257] ));
 sky130_fd_sc_hd__inv_2 \inv[1257]/_0_  (.A(\inv_in[1257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1258] ));
 sky130_fd_sc_hd__inv_2 \inv[1258]/_0_  (.A(\inv_in[1258] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1259] ));
 sky130_fd_sc_hd__inv_2 \inv[1259]/_0_  (.A(\inv_in[1259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1260] ));
 sky130_fd_sc_hd__inv_2 \inv[125]/_0_  (.A(\inv_in[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[126] ));
 sky130_fd_sc_hd__inv_2 \inv[1260]/_0_  (.A(\inv_in[1260] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1261] ));
 sky130_fd_sc_hd__inv_2 \inv[1261]/_0_  (.A(\inv_in[1261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1262] ));
 sky130_fd_sc_hd__inv_2 \inv[1262]/_0_  (.A(\inv_in[1262] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1263] ));
 sky130_fd_sc_hd__inv_2 \inv[1263]/_0_  (.A(\inv_in[1263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1264] ));
 sky130_fd_sc_hd__inv_2 \inv[1264]/_0_  (.A(\inv_in[1264] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1265] ));
 sky130_fd_sc_hd__inv_2 \inv[1265]/_0_  (.A(\inv_in[1265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1266] ));
 sky130_fd_sc_hd__inv_2 \inv[1266]/_0_  (.A(\inv_in[1266] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1267] ));
 sky130_fd_sc_hd__inv_2 \inv[1267]/_0_  (.A(\inv_in[1267] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1268] ));
 sky130_fd_sc_hd__inv_2 \inv[1268]/_0_  (.A(\inv_in[1268] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1269] ));
 sky130_fd_sc_hd__inv_2 \inv[1269]/_0_  (.A(\inv_in[1269] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1270] ));
 sky130_fd_sc_hd__inv_2 \inv[126]/_0_  (.A(\inv_in[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[127] ));
 sky130_fd_sc_hd__inv_2 \inv[1270]/_0_  (.A(\inv_in[1270] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1271] ));
 sky130_fd_sc_hd__inv_2 \inv[1271]/_0_  (.A(\inv_in[1271] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1272] ));
 sky130_fd_sc_hd__inv_2 \inv[1272]/_0_  (.A(\inv_in[1272] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1273] ));
 sky130_fd_sc_hd__inv_2 \inv[1273]/_0_  (.A(\inv_in[1273] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1274] ));
 sky130_fd_sc_hd__inv_2 \inv[1274]/_0_  (.A(\inv_in[1274] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1275] ));
 sky130_fd_sc_hd__inv_2 \inv[1275]/_0_  (.A(\inv_in[1275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1276] ));
 sky130_fd_sc_hd__inv_2 \inv[1276]/_0_  (.A(\inv_in[1276] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1277] ));
 sky130_fd_sc_hd__inv_2 \inv[1277]/_0_  (.A(\inv_in[1277] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1278] ));
 sky130_fd_sc_hd__inv_2 \inv[1278]/_0_  (.A(\inv_in[1278] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1279] ));
 sky130_fd_sc_hd__inv_2 \inv[1279]/_0_  (.A(\inv_in[1279] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1280] ));
 sky130_fd_sc_hd__inv_2 \inv[127]/_0_  (.A(\inv_in[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[128] ));
 sky130_fd_sc_hd__inv_2 \inv[1280]/_0_  (.A(\inv_in[1280] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1281] ));
 sky130_fd_sc_hd__inv_2 \inv[1281]/_0_  (.A(\inv_in[1281] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1282] ));
 sky130_fd_sc_hd__inv_2 \inv[1282]/_0_  (.A(\inv_in[1282] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1283] ));
 sky130_fd_sc_hd__inv_2 \inv[1283]/_0_  (.A(\inv_in[1283] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1284] ));
 sky130_fd_sc_hd__inv_2 \inv[1284]/_0_  (.A(\inv_in[1284] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1285] ));
 sky130_fd_sc_hd__inv_2 \inv[1285]/_0_  (.A(\inv_in[1285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1286] ));
 sky130_fd_sc_hd__inv_2 \inv[1286]/_0_  (.A(\inv_in[1286] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1287] ));
 sky130_fd_sc_hd__inv_2 \inv[1287]/_0_  (.A(\inv_in[1287] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1288] ));
 sky130_fd_sc_hd__inv_2 \inv[1288]/_0_  (.A(\inv_in[1288] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1289] ));
 sky130_fd_sc_hd__inv_2 \inv[1289]/_0_  (.A(\inv_in[1289] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1290] ));
 sky130_fd_sc_hd__inv_2 \inv[128]/_0_  (.A(\inv_in[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[129] ));
 sky130_fd_sc_hd__inv_2 \inv[1290]/_0_  (.A(\inv_in[1290] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1291] ));
 sky130_fd_sc_hd__inv_2 \inv[1291]/_0_  (.A(\inv_in[1291] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1292] ));
 sky130_fd_sc_hd__inv_2 \inv[1292]/_0_  (.A(\inv_in[1292] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1293] ));
 sky130_fd_sc_hd__inv_2 \inv[1293]/_0_  (.A(\inv_in[1293] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1294] ));
 sky130_fd_sc_hd__inv_2 \inv[1294]/_0_  (.A(\inv_in[1294] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1295] ));
 sky130_fd_sc_hd__inv_2 \inv[1295]/_0_  (.A(\inv_in[1295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1296] ));
 sky130_fd_sc_hd__inv_2 \inv[1296]/_0_  (.A(\inv_in[1296] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1297] ));
 sky130_fd_sc_hd__inv_2 \inv[1297]/_0_  (.A(\inv_in[1297] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1298] ));
 sky130_fd_sc_hd__inv_2 \inv[1298]/_0_  (.A(\inv_in[1298] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1299] ));
 sky130_fd_sc_hd__inv_2 \inv[1299]/_0_  (.A(\inv_in[1299] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1300] ));
 sky130_fd_sc_hd__inv_2 \inv[129]/_0_  (.A(\inv_in[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[130] ));
 sky130_fd_sc_hd__inv_2 \inv[12]/_0_  (.A(\inv_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[13] ));
 sky130_fd_sc_hd__inv_2 \inv[1300]/_0_  (.A(\inv_in[1300] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1301] ));
 sky130_fd_sc_hd__inv_2 \inv[1301]/_0_  (.A(\inv_in[1301] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1302] ));
 sky130_fd_sc_hd__inv_2 \inv[1302]/_0_  (.A(\inv_in[1302] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1303] ));
 sky130_fd_sc_hd__inv_2 \inv[1303]/_0_  (.A(\inv_in[1303] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1304] ));
 sky130_fd_sc_hd__inv_2 \inv[1304]/_0_  (.A(\inv_in[1304] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1305] ));
 sky130_fd_sc_hd__inv_2 \inv[1305]/_0_  (.A(\inv_in[1305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1306] ));
 sky130_fd_sc_hd__inv_2 \inv[1306]/_0_  (.A(\inv_in[1306] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1307] ));
 sky130_fd_sc_hd__inv_2 \inv[1307]/_0_  (.A(\inv_in[1307] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1308] ));
 sky130_fd_sc_hd__inv_2 \inv[1308]/_0_  (.A(\inv_in[1308] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1309] ));
 sky130_fd_sc_hd__inv_2 \inv[1309]/_0_  (.A(\inv_in[1309] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1310] ));
 sky130_fd_sc_hd__inv_2 \inv[130]/_0_  (.A(\inv_in[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[131] ));
 sky130_fd_sc_hd__inv_2 \inv[1310]/_0_  (.A(\inv_in[1310] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1311] ));
 sky130_fd_sc_hd__inv_2 \inv[1311]/_0_  (.A(\inv_in[1311] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1312] ));
 sky130_fd_sc_hd__inv_2 \inv[1312]/_0_  (.A(\inv_in[1312] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1313] ));
 sky130_fd_sc_hd__inv_2 \inv[1313]/_0_  (.A(\inv_in[1313] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1314] ));
 sky130_fd_sc_hd__inv_2 \inv[1314]/_0_  (.A(\inv_in[1314] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1315] ));
 sky130_fd_sc_hd__inv_2 \inv[1315]/_0_  (.A(\inv_in[1315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1316] ));
 sky130_fd_sc_hd__inv_2 \inv[1316]/_0_  (.A(\inv_in[1316] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1317] ));
 sky130_fd_sc_hd__inv_2 \inv[1317]/_0_  (.A(\inv_in[1317] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1318] ));
 sky130_fd_sc_hd__inv_2 \inv[1318]/_0_  (.A(\inv_in[1318] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1319] ));
 sky130_fd_sc_hd__inv_2 \inv[1319]/_0_  (.A(\inv_in[1319] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1320] ));
 sky130_fd_sc_hd__inv_2 \inv[131]/_0_  (.A(\inv_in[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[132] ));
 sky130_fd_sc_hd__inv_2 \inv[1320]/_0_  (.A(\inv_in[1320] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1321] ));
 sky130_fd_sc_hd__inv_2 \inv[1321]/_0_  (.A(\inv_in[1321] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1322] ));
 sky130_fd_sc_hd__inv_2 \inv[1322]/_0_  (.A(\inv_in[1322] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1323] ));
 sky130_fd_sc_hd__inv_2 \inv[1323]/_0_  (.A(\inv_in[1323] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1324] ));
 sky130_fd_sc_hd__inv_2 \inv[1324]/_0_  (.A(\inv_in[1324] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1325] ));
 sky130_fd_sc_hd__inv_2 \inv[1325]/_0_  (.A(\inv_in[1325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1326] ));
 sky130_fd_sc_hd__inv_2 \inv[1326]/_0_  (.A(\inv_in[1326] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1327] ));
 sky130_fd_sc_hd__inv_2 \inv[1327]/_0_  (.A(\inv_in[1327] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1328] ));
 sky130_fd_sc_hd__inv_2 \inv[1328]/_0_  (.A(\inv_in[1328] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1329] ));
 sky130_fd_sc_hd__inv_2 \inv[1329]/_0_  (.A(\inv_in[1329] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1330] ));
 sky130_fd_sc_hd__inv_2 \inv[132]/_0_  (.A(\inv_in[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[133] ));
 sky130_fd_sc_hd__inv_2 \inv[1330]/_0_  (.A(\inv_in[1330] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1331] ));
 sky130_fd_sc_hd__inv_2 \inv[1331]/_0_  (.A(\inv_in[1331] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1332] ));
 sky130_fd_sc_hd__inv_2 \inv[1332]/_0_  (.A(\inv_in[1332] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1333] ));
 sky130_fd_sc_hd__inv_2 \inv[1333]/_0_  (.A(\inv_in[1333] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1334] ));
 sky130_fd_sc_hd__inv_2 \inv[1334]/_0_  (.A(\inv_in[1334] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1335] ));
 sky130_fd_sc_hd__inv_2 \inv[1335]/_0_  (.A(\inv_in[1335] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1336] ));
 sky130_fd_sc_hd__inv_2 \inv[1336]/_0_  (.A(\inv_in[1336] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1337] ));
 sky130_fd_sc_hd__inv_2 \inv[1337]/_0_  (.A(\inv_in[1337] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1338] ));
 sky130_fd_sc_hd__inv_2 \inv[1338]/_0_  (.A(\inv_in[1338] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1339] ));
 sky130_fd_sc_hd__inv_2 \inv[1339]/_0_  (.A(\inv_in[1339] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1340] ));
 sky130_fd_sc_hd__inv_2 \inv[133]/_0_  (.A(\inv_in[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[134] ));
 sky130_fd_sc_hd__inv_2 \inv[1340]/_0_  (.A(\inv_in[1340] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1341] ));
 sky130_fd_sc_hd__inv_2 \inv[1341]/_0_  (.A(\inv_in[1341] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1342] ));
 sky130_fd_sc_hd__inv_2 \inv[1342]/_0_  (.A(\inv_in[1342] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1343] ));
 sky130_fd_sc_hd__inv_2 \inv[1343]/_0_  (.A(\inv_in[1343] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1344] ));
 sky130_fd_sc_hd__inv_2 \inv[1344]/_0_  (.A(\inv_in[1344] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1345] ));
 sky130_fd_sc_hd__inv_2 \inv[1345]/_0_  (.A(\inv_in[1345] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1346] ));
 sky130_fd_sc_hd__inv_2 \inv[1346]/_0_  (.A(\inv_in[1346] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1347] ));
 sky130_fd_sc_hd__inv_2 \inv[1347]/_0_  (.A(\inv_in[1347] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1348] ));
 sky130_fd_sc_hd__inv_2 \inv[1348]/_0_  (.A(\inv_in[1348] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1349] ));
 sky130_fd_sc_hd__inv_2 \inv[1349]/_0_  (.A(\inv_in[1349] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1350] ));
 sky130_fd_sc_hd__inv_2 \inv[134]/_0_  (.A(\inv_in[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[135] ));
 sky130_fd_sc_hd__inv_2 \inv[1350]/_0_  (.A(\inv_in[1350] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1351] ));
 sky130_fd_sc_hd__inv_2 \inv[1351]/_0_  (.A(\inv_in[1351] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1352] ));
 sky130_fd_sc_hd__inv_2 \inv[1352]/_0_  (.A(\inv_in[1352] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1353] ));
 sky130_fd_sc_hd__inv_2 \inv[1353]/_0_  (.A(\inv_in[1353] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1354] ));
 sky130_fd_sc_hd__inv_2 \inv[1354]/_0_  (.A(\inv_in[1354] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1355] ));
 sky130_fd_sc_hd__inv_2 \inv[1355]/_0_  (.A(\inv_in[1355] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1356] ));
 sky130_fd_sc_hd__inv_2 \inv[1356]/_0_  (.A(\inv_in[1356] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1357] ));
 sky130_fd_sc_hd__inv_2 \inv[1357]/_0_  (.A(\inv_in[1357] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1358] ));
 sky130_fd_sc_hd__inv_2 \inv[1358]/_0_  (.A(\inv_in[1358] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1359] ));
 sky130_fd_sc_hd__inv_2 \inv[1359]/_0_  (.A(\inv_in[1359] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1360] ));
 sky130_fd_sc_hd__inv_2 \inv[135]/_0_  (.A(\inv_in[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[136] ));
 sky130_fd_sc_hd__inv_2 \inv[1360]/_0_  (.A(\inv_in[1360] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1361] ));
 sky130_fd_sc_hd__inv_2 \inv[1361]/_0_  (.A(\inv_in[1361] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1362] ));
 sky130_fd_sc_hd__inv_2 \inv[1362]/_0_  (.A(\inv_in[1362] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1363] ));
 sky130_fd_sc_hd__inv_2 \inv[1363]/_0_  (.A(\inv_in[1363] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1364] ));
 sky130_fd_sc_hd__inv_2 \inv[1364]/_0_  (.A(\inv_in[1364] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1365] ));
 sky130_fd_sc_hd__inv_2 \inv[1365]/_0_  (.A(\inv_in[1365] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1366] ));
 sky130_fd_sc_hd__inv_2 \inv[1366]/_0_  (.A(\inv_in[1366] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1367] ));
 sky130_fd_sc_hd__inv_2 \inv[1367]/_0_  (.A(\inv_in[1367] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1368] ));
 sky130_fd_sc_hd__inv_2 \inv[1368]/_0_  (.A(\inv_in[1368] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1369] ));
 sky130_fd_sc_hd__inv_2 \inv[1369]/_0_  (.A(\inv_in[1369] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1370] ));
 sky130_fd_sc_hd__inv_2 \inv[136]/_0_  (.A(\inv_in[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[137] ));
 sky130_fd_sc_hd__inv_2 \inv[1370]/_0_  (.A(\inv_in[1370] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1371] ));
 sky130_fd_sc_hd__inv_2 \inv[1371]/_0_  (.A(\inv_in[1371] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1372] ));
 sky130_fd_sc_hd__inv_2 \inv[1372]/_0_  (.A(\inv_in[1372] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1373] ));
 sky130_fd_sc_hd__inv_2 \inv[1373]/_0_  (.A(\inv_in[1373] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1374] ));
 sky130_fd_sc_hd__inv_2 \inv[1374]/_0_  (.A(\inv_in[1374] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1375] ));
 sky130_fd_sc_hd__inv_2 \inv[1375]/_0_  (.A(\inv_in[1375] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1376] ));
 sky130_fd_sc_hd__inv_2 \inv[1376]/_0_  (.A(\inv_in[1376] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1377] ));
 sky130_fd_sc_hd__inv_2 \inv[1377]/_0_  (.A(\inv_in[1377] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1378] ));
 sky130_fd_sc_hd__inv_2 \inv[1378]/_0_  (.A(\inv_in[1378] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1379] ));
 sky130_fd_sc_hd__inv_2 \inv[1379]/_0_  (.A(\inv_in[1379] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1380] ));
 sky130_fd_sc_hd__inv_2 \inv[137]/_0_  (.A(\inv_in[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[138] ));
 sky130_fd_sc_hd__inv_2 \inv[1380]/_0_  (.A(\inv_in[1380] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1381] ));
 sky130_fd_sc_hd__inv_2 \inv[1381]/_0_  (.A(\inv_in[1381] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1382] ));
 sky130_fd_sc_hd__inv_2 \inv[1382]/_0_  (.A(\inv_in[1382] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1383] ));
 sky130_fd_sc_hd__inv_2 \inv[1383]/_0_  (.A(\inv_in[1383] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1384] ));
 sky130_fd_sc_hd__inv_2 \inv[1384]/_0_  (.A(\inv_in[1384] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1385] ));
 sky130_fd_sc_hd__inv_2 \inv[1385]/_0_  (.A(\inv_in[1385] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1386] ));
 sky130_fd_sc_hd__inv_2 \inv[1386]/_0_  (.A(\inv_in[1386] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1387] ));
 sky130_fd_sc_hd__inv_2 \inv[1387]/_0_  (.A(\inv_in[1387] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1388] ));
 sky130_fd_sc_hd__inv_2 \inv[1388]/_0_  (.A(\inv_in[1388] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1389] ));
 sky130_fd_sc_hd__inv_2 \inv[1389]/_0_  (.A(\inv_in[1389] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1390] ));
 sky130_fd_sc_hd__inv_2 \inv[138]/_0_  (.A(\inv_in[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[139] ));
 sky130_fd_sc_hd__inv_2 \inv[1390]/_0_  (.A(\inv_in[1390] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1391] ));
 sky130_fd_sc_hd__inv_2 \inv[1391]/_0_  (.A(\inv_in[1391] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1392] ));
 sky130_fd_sc_hd__inv_2 \inv[1392]/_0_  (.A(\inv_in[1392] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1393] ));
 sky130_fd_sc_hd__inv_2 \inv[1393]/_0_  (.A(\inv_in[1393] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1394] ));
 sky130_fd_sc_hd__inv_2 \inv[1394]/_0_  (.A(\inv_in[1394] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1395] ));
 sky130_fd_sc_hd__inv_2 \inv[1395]/_0_  (.A(\inv_in[1395] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1396] ));
 sky130_fd_sc_hd__inv_2 \inv[1396]/_0_  (.A(\inv_in[1396] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1397] ));
 sky130_fd_sc_hd__inv_2 \inv[1397]/_0_  (.A(\inv_in[1397] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1398] ));
 sky130_fd_sc_hd__inv_2 \inv[1398]/_0_  (.A(\inv_in[1398] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1399] ));
 sky130_fd_sc_hd__inv_2 \inv[1399]/_0_  (.A(\inv_in[1399] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1400] ));
 sky130_fd_sc_hd__inv_2 \inv[139]/_0_  (.A(\inv_in[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[140] ));
 sky130_fd_sc_hd__inv_2 \inv[13]/_0_  (.A(\inv_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[14] ));
 sky130_fd_sc_hd__inv_2 \inv[1400]/_0_  (.A(\inv_in[1400] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1401] ));
 sky130_fd_sc_hd__inv_2 \inv[1401]/_0_  (.A(\inv_in[1401] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1402] ));
 sky130_fd_sc_hd__inv_2 \inv[1402]/_0_  (.A(\inv_in[1402] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1403] ));
 sky130_fd_sc_hd__inv_2 \inv[1403]/_0_  (.A(\inv_in[1403] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1404] ));
 sky130_fd_sc_hd__inv_2 \inv[1404]/_0_  (.A(\inv_in[1404] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1405] ));
 sky130_fd_sc_hd__inv_2 \inv[1405]/_0_  (.A(\inv_in[1405] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1406] ));
 sky130_fd_sc_hd__inv_2 \inv[1406]/_0_  (.A(\inv_in[1406] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1407] ));
 sky130_fd_sc_hd__inv_2 \inv[1407]/_0_  (.A(\inv_in[1407] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1408] ));
 sky130_fd_sc_hd__inv_2 \inv[1408]/_0_  (.A(\inv_in[1408] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1409] ));
 sky130_fd_sc_hd__inv_2 \inv[1409]/_0_  (.A(\inv_in[1409] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1410] ));
 sky130_fd_sc_hd__inv_2 \inv[140]/_0_  (.A(\inv_in[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[141] ));
 sky130_fd_sc_hd__inv_2 \inv[1410]/_0_  (.A(\inv_in[1410] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1411] ));
 sky130_fd_sc_hd__inv_2 \inv[1411]/_0_  (.A(\inv_in[1411] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1412] ));
 sky130_fd_sc_hd__inv_2 \inv[1412]/_0_  (.A(\inv_in[1412] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1413] ));
 sky130_fd_sc_hd__inv_2 \inv[1413]/_0_  (.A(\inv_in[1413] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1414] ));
 sky130_fd_sc_hd__inv_2 \inv[1414]/_0_  (.A(\inv_in[1414] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1415] ));
 sky130_fd_sc_hd__inv_2 \inv[1415]/_0_  (.A(\inv_in[1415] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1416] ));
 sky130_fd_sc_hd__inv_2 \inv[1416]/_0_  (.A(\inv_in[1416] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1417] ));
 sky130_fd_sc_hd__inv_2 \inv[1417]/_0_  (.A(\inv_in[1417] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1418] ));
 sky130_fd_sc_hd__inv_2 \inv[1418]/_0_  (.A(\inv_in[1418] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1419] ));
 sky130_fd_sc_hd__inv_2 \inv[1419]/_0_  (.A(\inv_in[1419] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1420] ));
 sky130_fd_sc_hd__inv_2 \inv[141]/_0_  (.A(\inv_in[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[142] ));
 sky130_fd_sc_hd__inv_2 \inv[1420]/_0_  (.A(\inv_in[1420] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1421] ));
 sky130_fd_sc_hd__inv_2 \inv[1421]/_0_  (.A(\inv_in[1421] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1422] ));
 sky130_fd_sc_hd__inv_2 \inv[1422]/_0_  (.A(\inv_in[1422] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1423] ));
 sky130_fd_sc_hd__inv_2 \inv[1423]/_0_  (.A(\inv_in[1423] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1424] ));
 sky130_fd_sc_hd__inv_2 \inv[1424]/_0_  (.A(\inv_in[1424] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1425] ));
 sky130_fd_sc_hd__inv_2 \inv[1425]/_0_  (.A(\inv_in[1425] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1426] ));
 sky130_fd_sc_hd__inv_2 \inv[1426]/_0_  (.A(\inv_in[1426] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1427] ));
 sky130_fd_sc_hd__inv_2 \inv[1427]/_0_  (.A(\inv_in[1427] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1428] ));
 sky130_fd_sc_hd__inv_2 \inv[1428]/_0_  (.A(\inv_in[1428] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1429] ));
 sky130_fd_sc_hd__inv_2 \inv[1429]/_0_  (.A(\inv_in[1429] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1430] ));
 sky130_fd_sc_hd__inv_2 \inv[142]/_0_  (.A(\inv_in[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[143] ));
 sky130_fd_sc_hd__inv_2 \inv[1430]/_0_  (.A(\inv_in[1430] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1431] ));
 sky130_fd_sc_hd__inv_2 \inv[1431]/_0_  (.A(\inv_in[1431] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1432] ));
 sky130_fd_sc_hd__inv_2 \inv[1432]/_0_  (.A(\inv_in[1432] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1433] ));
 sky130_fd_sc_hd__inv_2 \inv[1433]/_0_  (.A(\inv_in[1433] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1434] ));
 sky130_fd_sc_hd__inv_2 \inv[1434]/_0_  (.A(\inv_in[1434] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1435] ));
 sky130_fd_sc_hd__inv_2 \inv[1435]/_0_  (.A(\inv_in[1435] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1436] ));
 sky130_fd_sc_hd__inv_2 \inv[1436]/_0_  (.A(\inv_in[1436] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1437] ));
 sky130_fd_sc_hd__inv_2 \inv[1437]/_0_  (.A(\inv_in[1437] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1438] ));
 sky130_fd_sc_hd__inv_2 \inv[1438]/_0_  (.A(\inv_in[1438] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1439] ));
 sky130_fd_sc_hd__inv_2 \inv[1439]/_0_  (.A(\inv_in[1439] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1440] ));
 sky130_fd_sc_hd__inv_2 \inv[143]/_0_  (.A(\inv_in[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[144] ));
 sky130_fd_sc_hd__inv_2 \inv[1440]/_0_  (.A(\inv_in[1440] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1441] ));
 sky130_fd_sc_hd__inv_2 \inv[1441]/_0_  (.A(\inv_in[1441] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1442] ));
 sky130_fd_sc_hd__inv_2 \inv[1442]/_0_  (.A(\inv_in[1442] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1443] ));
 sky130_fd_sc_hd__inv_2 \inv[1443]/_0_  (.A(\inv_in[1443] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1444] ));
 sky130_fd_sc_hd__inv_2 \inv[1444]/_0_  (.A(\inv_in[1444] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1445] ));
 sky130_fd_sc_hd__inv_2 \inv[1445]/_0_  (.A(\inv_in[1445] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1446] ));
 sky130_fd_sc_hd__inv_2 \inv[1446]/_0_  (.A(\inv_in[1446] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1447] ));
 sky130_fd_sc_hd__inv_2 \inv[1447]/_0_  (.A(\inv_in[1447] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1448] ));
 sky130_fd_sc_hd__inv_2 \inv[1448]/_0_  (.A(\inv_in[1448] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1449] ));
 sky130_fd_sc_hd__inv_2 \inv[1449]/_0_  (.A(\inv_in[1449] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1450] ));
 sky130_fd_sc_hd__inv_2 \inv[144]/_0_  (.A(\inv_in[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[145] ));
 sky130_fd_sc_hd__inv_2 \inv[1450]/_0_  (.A(\inv_in[1450] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1451] ));
 sky130_fd_sc_hd__inv_2 \inv[1451]/_0_  (.A(\inv_in[1451] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1452] ));
 sky130_fd_sc_hd__inv_2 \inv[1452]/_0_  (.A(\inv_in[1452] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1453] ));
 sky130_fd_sc_hd__inv_2 \inv[1453]/_0_  (.A(\inv_in[1453] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1454] ));
 sky130_fd_sc_hd__inv_2 \inv[1454]/_0_  (.A(\inv_in[1454] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1455] ));
 sky130_fd_sc_hd__inv_2 \inv[1455]/_0_  (.A(\inv_in[1455] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1456] ));
 sky130_fd_sc_hd__inv_2 \inv[1456]/_0_  (.A(\inv_in[1456] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1457] ));
 sky130_fd_sc_hd__inv_2 \inv[1457]/_0_  (.A(\inv_in[1457] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1458] ));
 sky130_fd_sc_hd__inv_2 \inv[1458]/_0_  (.A(\inv_in[1458] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1459] ));
 sky130_fd_sc_hd__inv_2 \inv[1459]/_0_  (.A(\inv_in[1459] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1460] ));
 sky130_fd_sc_hd__inv_2 \inv[145]/_0_  (.A(\inv_in[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[146] ));
 sky130_fd_sc_hd__inv_2 \inv[1460]/_0_  (.A(\inv_in[1460] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1461] ));
 sky130_fd_sc_hd__inv_2 \inv[1461]/_0_  (.A(\inv_in[1461] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1462] ));
 sky130_fd_sc_hd__inv_2 \inv[1462]/_0_  (.A(\inv_in[1462] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1463] ));
 sky130_fd_sc_hd__inv_2 \inv[1463]/_0_  (.A(\inv_in[1463] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1464] ));
 sky130_fd_sc_hd__inv_2 \inv[1464]/_0_  (.A(\inv_in[1464] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1465] ));
 sky130_fd_sc_hd__inv_2 \inv[1465]/_0_  (.A(\inv_in[1465] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1466] ));
 sky130_fd_sc_hd__inv_2 \inv[1466]/_0_  (.A(\inv_in[1466] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1467] ));
 sky130_fd_sc_hd__inv_2 \inv[1467]/_0_  (.A(\inv_in[1467] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1468] ));
 sky130_fd_sc_hd__inv_2 \inv[1468]/_0_  (.A(\inv_in[1468] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1469] ));
 sky130_fd_sc_hd__inv_2 \inv[1469]/_0_  (.A(\inv_in[1469] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1470] ));
 sky130_fd_sc_hd__inv_2 \inv[146]/_0_  (.A(\inv_in[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[147] ));
 sky130_fd_sc_hd__inv_2 \inv[1470]/_0_  (.A(\inv_in[1470] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1471] ));
 sky130_fd_sc_hd__inv_2 \inv[1471]/_0_  (.A(\inv_in[1471] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1472] ));
 sky130_fd_sc_hd__inv_2 \inv[1472]/_0_  (.A(\inv_in[1472] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1473] ));
 sky130_fd_sc_hd__inv_2 \inv[1473]/_0_  (.A(\inv_in[1473] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1474] ));
 sky130_fd_sc_hd__inv_2 \inv[1474]/_0_  (.A(\inv_in[1474] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1475] ));
 sky130_fd_sc_hd__inv_2 \inv[1475]/_0_  (.A(\inv_in[1475] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1476] ));
 sky130_fd_sc_hd__inv_2 \inv[1476]/_0_  (.A(\inv_in[1476] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1477] ));
 sky130_fd_sc_hd__inv_2 \inv[1477]/_0_  (.A(\inv_in[1477] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1478] ));
 sky130_fd_sc_hd__inv_2 \inv[1478]/_0_  (.A(\inv_in[1478] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1479] ));
 sky130_fd_sc_hd__inv_2 \inv[1479]/_0_  (.A(\inv_in[1479] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1480] ));
 sky130_fd_sc_hd__inv_2 \inv[147]/_0_  (.A(\inv_in[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[148] ));
 sky130_fd_sc_hd__inv_2 \inv[1480]/_0_  (.A(\inv_in[1480] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1481] ));
 sky130_fd_sc_hd__inv_2 \inv[1481]/_0_  (.A(\inv_in[1481] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1482] ));
 sky130_fd_sc_hd__inv_2 \inv[1482]/_0_  (.A(\inv_in[1482] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1483] ));
 sky130_fd_sc_hd__inv_2 \inv[1483]/_0_  (.A(\inv_in[1483] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1484] ));
 sky130_fd_sc_hd__inv_2 \inv[1484]/_0_  (.A(\inv_in[1484] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1485] ));
 sky130_fd_sc_hd__inv_2 \inv[1485]/_0_  (.A(\inv_in[1485] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1486] ));
 sky130_fd_sc_hd__inv_2 \inv[1486]/_0_  (.A(\inv_in[1486] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1487] ));
 sky130_fd_sc_hd__inv_2 \inv[1487]/_0_  (.A(\inv_in[1487] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1488] ));
 sky130_fd_sc_hd__inv_2 \inv[1488]/_0_  (.A(\inv_in[1488] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1489] ));
 sky130_fd_sc_hd__inv_2 \inv[1489]/_0_  (.A(\inv_in[1489] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1490] ));
 sky130_fd_sc_hd__inv_2 \inv[148]/_0_  (.A(\inv_in[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[149] ));
 sky130_fd_sc_hd__inv_2 \inv[1490]/_0_  (.A(\inv_in[1490] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1491] ));
 sky130_fd_sc_hd__inv_2 \inv[1491]/_0_  (.A(\inv_in[1491] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1492] ));
 sky130_fd_sc_hd__inv_2 \inv[1492]/_0_  (.A(\inv_in[1492] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1493] ));
 sky130_fd_sc_hd__inv_2 \inv[1493]/_0_  (.A(\inv_in[1493] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1494] ));
 sky130_fd_sc_hd__inv_2 \inv[1494]/_0_  (.A(\inv_in[1494] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1495] ));
 sky130_fd_sc_hd__inv_2 \inv[1495]/_0_  (.A(\inv_in[1495] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1496] ));
 sky130_fd_sc_hd__inv_2 \inv[1496]/_0_  (.A(\inv_in[1496] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1497] ));
 sky130_fd_sc_hd__inv_2 \inv[1497]/_0_  (.A(\inv_in[1497] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1498] ));
 sky130_fd_sc_hd__inv_2 \inv[1498]/_0_  (.A(\inv_in[1498] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1499] ));
 sky130_fd_sc_hd__inv_2 \inv[1499]/_0_  (.A(\inv_in[1499] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1500] ));
 sky130_fd_sc_hd__inv_2 \inv[149]/_0_  (.A(\inv_in[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[150] ));
 sky130_fd_sc_hd__inv_2 \inv[14]/_0_  (.A(\inv_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[15] ));
 sky130_fd_sc_hd__inv_2 \inv[1500]/_0_  (.A(\inv_in[1500] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1501] ));
 sky130_fd_sc_hd__inv_2 \inv[1501]/_0_  (.A(\inv_in[1501] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1502] ));
 sky130_fd_sc_hd__inv_2 \inv[1502]/_0_  (.A(\inv_in[1502] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1503] ));
 sky130_fd_sc_hd__inv_2 \inv[1503]/_0_  (.A(\inv_in[1503] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1504] ));
 sky130_fd_sc_hd__inv_2 \inv[1504]/_0_  (.A(\inv_in[1504] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1505] ));
 sky130_fd_sc_hd__inv_2 \inv[1505]/_0_  (.A(\inv_in[1505] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1506] ));
 sky130_fd_sc_hd__inv_2 \inv[1506]/_0_  (.A(\inv_in[1506] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1507] ));
 sky130_fd_sc_hd__inv_2 \inv[1507]/_0_  (.A(\inv_in[1507] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1508] ));
 sky130_fd_sc_hd__inv_2 \inv[1508]/_0_  (.A(\inv_in[1508] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1509] ));
 sky130_fd_sc_hd__inv_2 \inv[1509]/_0_  (.A(\inv_in[1509] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1510] ));
 sky130_fd_sc_hd__inv_2 \inv[150]/_0_  (.A(\inv_in[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[151] ));
 sky130_fd_sc_hd__inv_2 \inv[1510]/_0_  (.A(\inv_in[1510] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1511] ));
 sky130_fd_sc_hd__inv_2 \inv[1511]/_0_  (.A(\inv_in[1511] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1512] ));
 sky130_fd_sc_hd__inv_2 \inv[1512]/_0_  (.A(\inv_in[1512] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1513] ));
 sky130_fd_sc_hd__inv_2 \inv[1513]/_0_  (.A(\inv_in[1513] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1514] ));
 sky130_fd_sc_hd__inv_2 \inv[1514]/_0_  (.A(\inv_in[1514] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1515] ));
 sky130_fd_sc_hd__inv_2 \inv[1515]/_0_  (.A(\inv_in[1515] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1516] ));
 sky130_fd_sc_hd__inv_2 \inv[1516]/_0_  (.A(\inv_in[1516] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1517] ));
 sky130_fd_sc_hd__inv_2 \inv[1517]/_0_  (.A(\inv_in[1517] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1518] ));
 sky130_fd_sc_hd__inv_2 \inv[1518]/_0_  (.A(\inv_in[1518] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1519] ));
 sky130_fd_sc_hd__inv_2 \inv[1519]/_0_  (.A(\inv_in[1519] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1520] ));
 sky130_fd_sc_hd__inv_2 \inv[151]/_0_  (.A(\inv_in[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[152] ));
 sky130_fd_sc_hd__inv_2 \inv[1520]/_0_  (.A(\inv_in[1520] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1521] ));
 sky130_fd_sc_hd__inv_2 \inv[1521]/_0_  (.A(\inv_in[1521] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1522] ));
 sky130_fd_sc_hd__inv_2 \inv[1522]/_0_  (.A(\inv_in[1522] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1523] ));
 sky130_fd_sc_hd__inv_2 \inv[1523]/_0_  (.A(\inv_in[1523] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1524] ));
 sky130_fd_sc_hd__inv_2 \inv[1524]/_0_  (.A(\inv_in[1524] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1525] ));
 sky130_fd_sc_hd__inv_2 \inv[1525]/_0_  (.A(\inv_in[1525] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1526] ));
 sky130_fd_sc_hd__inv_2 \inv[1526]/_0_  (.A(\inv_in[1526] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1527] ));
 sky130_fd_sc_hd__inv_2 \inv[1527]/_0_  (.A(\inv_in[1527] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1528] ));
 sky130_fd_sc_hd__inv_2 \inv[1528]/_0_  (.A(\inv_in[1528] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1529] ));
 sky130_fd_sc_hd__inv_2 \inv[1529]/_0_  (.A(\inv_in[1529] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1530] ));
 sky130_fd_sc_hd__inv_2 \inv[152]/_0_  (.A(\inv_in[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[153] ));
 sky130_fd_sc_hd__inv_2 \inv[1530]/_0_  (.A(\inv_in[1530] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1531] ));
 sky130_fd_sc_hd__inv_2 \inv[1531]/_0_  (.A(\inv_in[1531] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1532] ));
 sky130_fd_sc_hd__inv_2 \inv[1532]/_0_  (.A(\inv_in[1532] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1533] ));
 sky130_fd_sc_hd__inv_2 \inv[1533]/_0_  (.A(\inv_in[1533] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1534] ));
 sky130_fd_sc_hd__inv_2 \inv[1534]/_0_  (.A(\inv_in[1534] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1535] ));
 sky130_fd_sc_hd__inv_2 \inv[1535]/_0_  (.A(\inv_in[1535] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1536] ));
 sky130_fd_sc_hd__inv_2 \inv[1536]/_0_  (.A(\inv_in[1536] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1537] ));
 sky130_fd_sc_hd__inv_2 \inv[1537]/_0_  (.A(\inv_in[1537] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1538] ));
 sky130_fd_sc_hd__inv_2 \inv[1538]/_0_  (.A(\inv_in[1538] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1539] ));
 sky130_fd_sc_hd__inv_2 \inv[1539]/_0_  (.A(\inv_in[1539] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1540] ));
 sky130_fd_sc_hd__inv_2 \inv[153]/_0_  (.A(\inv_in[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[154] ));
 sky130_fd_sc_hd__inv_2 \inv[1540]/_0_  (.A(\inv_in[1540] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1541] ));
 sky130_fd_sc_hd__inv_2 \inv[1541]/_0_  (.A(\inv_in[1541] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1542] ));
 sky130_fd_sc_hd__inv_2 \inv[1542]/_0_  (.A(\inv_in[1542] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1543] ));
 sky130_fd_sc_hd__inv_2 \inv[1543]/_0_  (.A(\inv_in[1543] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1544] ));
 sky130_fd_sc_hd__inv_2 \inv[1544]/_0_  (.A(\inv_in[1544] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1545] ));
 sky130_fd_sc_hd__inv_2 \inv[1545]/_0_  (.A(\inv_in[1545] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1546] ));
 sky130_fd_sc_hd__inv_2 \inv[1546]/_0_  (.A(\inv_in[1546] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1547] ));
 sky130_fd_sc_hd__inv_2 \inv[1547]/_0_  (.A(\inv_in[1547] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1548] ));
 sky130_fd_sc_hd__inv_2 \inv[1548]/_0_  (.A(\inv_in[1548] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1549] ));
 sky130_fd_sc_hd__inv_2 \inv[1549]/_0_  (.A(\inv_in[1549] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1550] ));
 sky130_fd_sc_hd__inv_2 \inv[154]/_0_  (.A(\inv_in[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[155] ));
 sky130_fd_sc_hd__inv_2 \inv[1550]/_0_  (.A(\inv_in[1550] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1551] ));
 sky130_fd_sc_hd__inv_2 \inv[1551]/_0_  (.A(\inv_in[1551] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1552] ));
 sky130_fd_sc_hd__inv_2 \inv[1552]/_0_  (.A(\inv_in[1552] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1553] ));
 sky130_fd_sc_hd__inv_2 \inv[1553]/_0_  (.A(\inv_in[1553] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1554] ));
 sky130_fd_sc_hd__inv_2 \inv[1554]/_0_  (.A(\inv_in[1554] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1555] ));
 sky130_fd_sc_hd__inv_2 \inv[1555]/_0_  (.A(\inv_in[1555] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1556] ));
 sky130_fd_sc_hd__inv_2 \inv[1556]/_0_  (.A(\inv_in[1556] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1557] ));
 sky130_fd_sc_hd__inv_2 \inv[1557]/_0_  (.A(\inv_in[1557] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1558] ));
 sky130_fd_sc_hd__inv_2 \inv[1558]/_0_  (.A(\inv_in[1558] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1559] ));
 sky130_fd_sc_hd__inv_2 \inv[1559]/_0_  (.A(\inv_in[1559] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1560] ));
 sky130_fd_sc_hd__inv_2 \inv[155]/_0_  (.A(\inv_in[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[156] ));
 sky130_fd_sc_hd__inv_2 \inv[1560]/_0_  (.A(\inv_in[1560] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1561] ));
 sky130_fd_sc_hd__inv_2 \inv[1561]/_0_  (.A(\inv_in[1561] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1562] ));
 sky130_fd_sc_hd__inv_2 \inv[1562]/_0_  (.A(\inv_in[1562] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1563] ));
 sky130_fd_sc_hd__inv_2 \inv[1563]/_0_  (.A(\inv_in[1563] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1564] ));
 sky130_fd_sc_hd__inv_2 \inv[1564]/_0_  (.A(\inv_in[1564] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1565] ));
 sky130_fd_sc_hd__inv_2 \inv[1565]/_0_  (.A(\inv_in[1565] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1566] ));
 sky130_fd_sc_hd__inv_2 \inv[1566]/_0_  (.A(\inv_in[1566] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1567] ));
 sky130_fd_sc_hd__inv_2 \inv[1567]/_0_  (.A(\inv_in[1567] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1568] ));
 sky130_fd_sc_hd__inv_2 \inv[1568]/_0_  (.A(\inv_in[1568] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1569] ));
 sky130_fd_sc_hd__inv_2 \inv[1569]/_0_  (.A(\inv_in[1569] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1570] ));
 sky130_fd_sc_hd__inv_2 \inv[156]/_0_  (.A(\inv_in[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[157] ));
 sky130_fd_sc_hd__inv_2 \inv[1570]/_0_  (.A(\inv_in[1570] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1571] ));
 sky130_fd_sc_hd__inv_2 \inv[1571]/_0_  (.A(\inv_in[1571] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1572] ));
 sky130_fd_sc_hd__inv_2 \inv[1572]/_0_  (.A(\inv_in[1572] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1573] ));
 sky130_fd_sc_hd__inv_2 \inv[1573]/_0_  (.A(\inv_in[1573] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1574] ));
 sky130_fd_sc_hd__inv_2 \inv[1574]/_0_  (.A(\inv_in[1574] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1575] ));
 sky130_fd_sc_hd__inv_2 \inv[1575]/_0_  (.A(\inv_in[1575] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1576] ));
 sky130_fd_sc_hd__inv_2 \inv[1576]/_0_  (.A(\inv_in[1576] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1577] ));
 sky130_fd_sc_hd__inv_2 \inv[1577]/_0_  (.A(\inv_in[1577] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1578] ));
 sky130_fd_sc_hd__inv_2 \inv[1578]/_0_  (.A(\inv_in[1578] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1579] ));
 sky130_fd_sc_hd__inv_2 \inv[1579]/_0_  (.A(\inv_in[1579] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1580] ));
 sky130_fd_sc_hd__inv_2 \inv[157]/_0_  (.A(\inv_in[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[158] ));
 sky130_fd_sc_hd__inv_2 \inv[1580]/_0_  (.A(\inv_in[1580] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1581] ));
 sky130_fd_sc_hd__inv_2 \inv[1581]/_0_  (.A(\inv_in[1581] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1582] ));
 sky130_fd_sc_hd__inv_2 \inv[1582]/_0_  (.A(\inv_in[1582] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1583] ));
 sky130_fd_sc_hd__inv_2 \inv[1583]/_0_  (.A(\inv_in[1583] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1584] ));
 sky130_fd_sc_hd__inv_2 \inv[1584]/_0_  (.A(\inv_in[1584] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1585] ));
 sky130_fd_sc_hd__inv_2 \inv[1585]/_0_  (.A(\inv_in[1585] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1586] ));
 sky130_fd_sc_hd__inv_2 \inv[1586]/_0_  (.A(\inv_in[1586] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1587] ));
 sky130_fd_sc_hd__inv_2 \inv[1587]/_0_  (.A(\inv_in[1587] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1588] ));
 sky130_fd_sc_hd__inv_2 \inv[1588]/_0_  (.A(\inv_in[1588] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1589] ));
 sky130_fd_sc_hd__inv_2 \inv[1589]/_0_  (.A(\inv_in[1589] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1590] ));
 sky130_fd_sc_hd__inv_2 \inv[158]/_0_  (.A(\inv_in[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[159] ));
 sky130_fd_sc_hd__inv_2 \inv[1590]/_0_  (.A(\inv_in[1590] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1591] ));
 sky130_fd_sc_hd__inv_2 \inv[1591]/_0_  (.A(\inv_in[1591] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1592] ));
 sky130_fd_sc_hd__inv_2 \inv[1592]/_0_  (.A(\inv_in[1592] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1593] ));
 sky130_fd_sc_hd__inv_2 \inv[1593]/_0_  (.A(\inv_in[1593] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1594] ));
 sky130_fd_sc_hd__inv_2 \inv[1594]/_0_  (.A(\inv_in[1594] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1595] ));
 sky130_fd_sc_hd__inv_2 \inv[1595]/_0_  (.A(\inv_in[1595] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1596] ));
 sky130_fd_sc_hd__inv_2 \inv[1596]/_0_  (.A(\inv_in[1596] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1597] ));
 sky130_fd_sc_hd__inv_2 \inv[1597]/_0_  (.A(\inv_in[1597] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1598] ));
 sky130_fd_sc_hd__inv_2 \inv[1598]/_0_  (.A(\inv_in[1598] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1599] ));
 sky130_fd_sc_hd__inv_2 \inv[1599]/_0_  (.A(\inv_in[1599] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1600] ));
 sky130_fd_sc_hd__inv_2 \inv[159]/_0_  (.A(\inv_in[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[160] ));
 sky130_fd_sc_hd__inv_2 \inv[15]/_0_  (.A(\inv_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[16] ));
 sky130_fd_sc_hd__inv_2 \inv[1600]/_0_  (.A(\inv_in[1600] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1601] ));
 sky130_fd_sc_hd__inv_2 \inv[1601]/_0_  (.A(\inv_in[1601] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1602] ));
 sky130_fd_sc_hd__inv_2 \inv[1602]/_0_  (.A(\inv_in[1602] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1603] ));
 sky130_fd_sc_hd__inv_2 \inv[1603]/_0_  (.A(\inv_in[1603] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1604] ));
 sky130_fd_sc_hd__inv_2 \inv[1604]/_0_  (.A(\inv_in[1604] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1605] ));
 sky130_fd_sc_hd__inv_2 \inv[1605]/_0_  (.A(\inv_in[1605] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1606] ));
 sky130_fd_sc_hd__inv_2 \inv[1606]/_0_  (.A(\inv_in[1606] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1607] ));
 sky130_fd_sc_hd__inv_2 \inv[1607]/_0_  (.A(\inv_in[1607] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1608] ));
 sky130_fd_sc_hd__inv_2 \inv[1608]/_0_  (.A(\inv_in[1608] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1609] ));
 sky130_fd_sc_hd__inv_2 \inv[1609]/_0_  (.A(\inv_in[1609] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1610] ));
 sky130_fd_sc_hd__inv_2 \inv[160]/_0_  (.A(\inv_in[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[161] ));
 sky130_fd_sc_hd__inv_2 \inv[1610]/_0_  (.A(\inv_in[1610] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1611] ));
 sky130_fd_sc_hd__inv_2 \inv[1611]/_0_  (.A(\inv_in[1611] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1612] ));
 sky130_fd_sc_hd__inv_2 \inv[1612]/_0_  (.A(\inv_in[1612] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1613] ));
 sky130_fd_sc_hd__inv_2 \inv[1613]/_0_  (.A(\inv_in[1613] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1614] ));
 sky130_fd_sc_hd__inv_2 \inv[1614]/_0_  (.A(\inv_in[1614] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1615] ));
 sky130_fd_sc_hd__inv_2 \inv[1615]/_0_  (.A(\inv_in[1615] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1616] ));
 sky130_fd_sc_hd__inv_2 \inv[1616]/_0_  (.A(\inv_in[1616] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1617] ));
 sky130_fd_sc_hd__inv_2 \inv[1617]/_0_  (.A(\inv_in[1617] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1618] ));
 sky130_fd_sc_hd__inv_2 \inv[1618]/_0_  (.A(\inv_in[1618] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1619] ));
 sky130_fd_sc_hd__inv_2 \inv[1619]/_0_  (.A(\inv_in[1619] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1620] ));
 sky130_fd_sc_hd__inv_2 \inv[161]/_0_  (.A(\inv_in[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[162] ));
 sky130_fd_sc_hd__inv_2 \inv[1620]/_0_  (.A(\inv_in[1620] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1621] ));
 sky130_fd_sc_hd__inv_2 \inv[1621]/_0_  (.A(\inv_in[1621] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1622] ));
 sky130_fd_sc_hd__inv_2 \inv[1622]/_0_  (.A(\inv_in[1622] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1623] ));
 sky130_fd_sc_hd__inv_2 \inv[1623]/_0_  (.A(\inv_in[1623] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1624] ));
 sky130_fd_sc_hd__inv_2 \inv[1624]/_0_  (.A(\inv_in[1624] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1625] ));
 sky130_fd_sc_hd__inv_2 \inv[1625]/_0_  (.A(\inv_in[1625] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1626] ));
 sky130_fd_sc_hd__inv_2 \inv[1626]/_0_  (.A(\inv_in[1626] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1627] ));
 sky130_fd_sc_hd__inv_2 \inv[1627]/_0_  (.A(\inv_in[1627] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1628] ));
 sky130_fd_sc_hd__inv_2 \inv[1628]/_0_  (.A(\inv_in[1628] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1629] ));
 sky130_fd_sc_hd__inv_2 \inv[1629]/_0_  (.A(\inv_in[1629] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1630] ));
 sky130_fd_sc_hd__inv_2 \inv[162]/_0_  (.A(\inv_in[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[163] ));
 sky130_fd_sc_hd__inv_2 \inv[1630]/_0_  (.A(\inv_in[1630] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1631] ));
 sky130_fd_sc_hd__inv_2 \inv[1631]/_0_  (.A(\inv_in[1631] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1632] ));
 sky130_fd_sc_hd__inv_2 \inv[1632]/_0_  (.A(\inv_in[1632] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1633] ));
 sky130_fd_sc_hd__inv_2 \inv[1633]/_0_  (.A(\inv_in[1633] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1634] ));
 sky130_fd_sc_hd__inv_2 \inv[1634]/_0_  (.A(\inv_in[1634] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1635] ));
 sky130_fd_sc_hd__inv_2 \inv[1635]/_0_  (.A(\inv_in[1635] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1636] ));
 sky130_fd_sc_hd__inv_2 \inv[1636]/_0_  (.A(\inv_in[1636] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1637] ));
 sky130_fd_sc_hd__inv_2 \inv[1637]/_0_  (.A(\inv_in[1637] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1638] ));
 sky130_fd_sc_hd__inv_2 \inv[1638]/_0_  (.A(\inv_in[1638] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1639] ));
 sky130_fd_sc_hd__inv_2 \inv[1639]/_0_  (.A(\inv_in[1639] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1640] ));
 sky130_fd_sc_hd__inv_2 \inv[163]/_0_  (.A(\inv_in[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[164] ));
 sky130_fd_sc_hd__inv_2 \inv[1640]/_0_  (.A(\inv_in[1640] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1641] ));
 sky130_fd_sc_hd__inv_2 \inv[1641]/_0_  (.A(\inv_in[1641] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1642] ));
 sky130_fd_sc_hd__inv_2 \inv[1642]/_0_  (.A(\inv_in[1642] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1643] ));
 sky130_fd_sc_hd__inv_2 \inv[1643]/_0_  (.A(\inv_in[1643] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1644] ));
 sky130_fd_sc_hd__inv_2 \inv[1644]/_0_  (.A(\inv_in[1644] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1645] ));
 sky130_fd_sc_hd__inv_2 \inv[1645]/_0_  (.A(\inv_in[1645] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1646] ));
 sky130_fd_sc_hd__inv_2 \inv[1646]/_0_  (.A(\inv_in[1646] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1647] ));
 sky130_fd_sc_hd__inv_2 \inv[1647]/_0_  (.A(\inv_in[1647] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1648] ));
 sky130_fd_sc_hd__inv_2 \inv[1648]/_0_  (.A(\inv_in[1648] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1649] ));
 sky130_fd_sc_hd__inv_2 \inv[1649]/_0_  (.A(\inv_in[1649] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1650] ));
 sky130_fd_sc_hd__inv_2 \inv[164]/_0_  (.A(\inv_in[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[165] ));
 sky130_fd_sc_hd__inv_2 \inv[1650]/_0_  (.A(\inv_in[1650] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1651] ));
 sky130_fd_sc_hd__inv_2 \inv[1651]/_0_  (.A(\inv_in[1651] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1652] ));
 sky130_fd_sc_hd__inv_2 \inv[1652]/_0_  (.A(\inv_in[1652] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1653] ));
 sky130_fd_sc_hd__inv_2 \inv[1653]/_0_  (.A(\inv_in[1653] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1654] ));
 sky130_fd_sc_hd__inv_2 \inv[1654]/_0_  (.A(\inv_in[1654] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1655] ));
 sky130_fd_sc_hd__inv_2 \inv[1655]/_0_  (.A(\inv_in[1655] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1656] ));
 sky130_fd_sc_hd__inv_2 \inv[1656]/_0_  (.A(\inv_in[1656] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1657] ));
 sky130_fd_sc_hd__inv_2 \inv[1657]/_0_  (.A(\inv_in[1657] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1658] ));
 sky130_fd_sc_hd__inv_2 \inv[1658]/_0_  (.A(\inv_in[1658] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1659] ));
 sky130_fd_sc_hd__inv_2 \inv[1659]/_0_  (.A(\inv_in[1659] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1660] ));
 sky130_fd_sc_hd__inv_2 \inv[165]/_0_  (.A(\inv_in[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[166] ));
 sky130_fd_sc_hd__inv_2 \inv[1660]/_0_  (.A(\inv_in[1660] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1661] ));
 sky130_fd_sc_hd__inv_2 \inv[1661]/_0_  (.A(\inv_in[1661] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1662] ));
 sky130_fd_sc_hd__inv_2 \inv[1662]/_0_  (.A(\inv_in[1662] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1663] ));
 sky130_fd_sc_hd__inv_2 \inv[1663]/_0_  (.A(\inv_in[1663] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1664] ));
 sky130_fd_sc_hd__inv_2 \inv[1664]/_0_  (.A(\inv_in[1664] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1665] ));
 sky130_fd_sc_hd__inv_2 \inv[1665]/_0_  (.A(\inv_in[1665] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1666] ));
 sky130_fd_sc_hd__inv_2 \inv[1666]/_0_  (.A(\inv_in[1666] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1667] ));
 sky130_fd_sc_hd__inv_2 \inv[1667]/_0_  (.A(\inv_in[1667] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1668] ));
 sky130_fd_sc_hd__inv_2 \inv[1668]/_0_  (.A(\inv_in[1668] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1669] ));
 sky130_fd_sc_hd__inv_2 \inv[1669]/_0_  (.A(\inv_in[1669] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1670] ));
 sky130_fd_sc_hd__inv_2 \inv[166]/_0_  (.A(\inv_in[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[167] ));
 sky130_fd_sc_hd__inv_2 \inv[1670]/_0_  (.A(\inv_in[1670] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1671] ));
 sky130_fd_sc_hd__inv_2 \inv[1671]/_0_  (.A(\inv_in[1671] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1672] ));
 sky130_fd_sc_hd__inv_2 \inv[1672]/_0_  (.A(\inv_in[1672] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1673] ));
 sky130_fd_sc_hd__inv_2 \inv[1673]/_0_  (.A(\inv_in[1673] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1674] ));
 sky130_fd_sc_hd__inv_2 \inv[1674]/_0_  (.A(\inv_in[1674] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1675] ));
 sky130_fd_sc_hd__inv_2 \inv[1675]/_0_  (.A(\inv_in[1675] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1676] ));
 sky130_fd_sc_hd__inv_2 \inv[1676]/_0_  (.A(\inv_in[1676] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1677] ));
 sky130_fd_sc_hd__inv_2 \inv[1677]/_0_  (.A(\inv_in[1677] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1678] ));
 sky130_fd_sc_hd__inv_2 \inv[1678]/_0_  (.A(\inv_in[1678] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1679] ));
 sky130_fd_sc_hd__inv_2 \inv[1679]/_0_  (.A(\inv_in[1679] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1680] ));
 sky130_fd_sc_hd__inv_2 \inv[167]/_0_  (.A(\inv_in[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[168] ));
 sky130_fd_sc_hd__inv_2 \inv[1680]/_0_  (.A(\inv_in[1680] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1681] ));
 sky130_fd_sc_hd__inv_2 \inv[1681]/_0_  (.A(\inv_in[1681] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1682] ));
 sky130_fd_sc_hd__inv_2 \inv[1682]/_0_  (.A(\inv_in[1682] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1683] ));
 sky130_fd_sc_hd__inv_2 \inv[1683]/_0_  (.A(\inv_in[1683] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1684] ));
 sky130_fd_sc_hd__inv_2 \inv[1684]/_0_  (.A(\inv_in[1684] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1685] ));
 sky130_fd_sc_hd__inv_2 \inv[1685]/_0_  (.A(\inv_in[1685] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1686] ));
 sky130_fd_sc_hd__inv_2 \inv[1686]/_0_  (.A(\inv_in[1686] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1687] ));
 sky130_fd_sc_hd__inv_2 \inv[1687]/_0_  (.A(\inv_in[1687] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1688] ));
 sky130_fd_sc_hd__inv_2 \inv[1688]/_0_  (.A(\inv_in[1688] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1689] ));
 sky130_fd_sc_hd__inv_2 \inv[1689]/_0_  (.A(\inv_in[1689] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1690] ));
 sky130_fd_sc_hd__inv_2 \inv[168]/_0_  (.A(\inv_in[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[169] ));
 sky130_fd_sc_hd__inv_2 \inv[1690]/_0_  (.A(\inv_in[1690] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1691] ));
 sky130_fd_sc_hd__inv_2 \inv[1691]/_0_  (.A(\inv_in[1691] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1692] ));
 sky130_fd_sc_hd__inv_2 \inv[1692]/_0_  (.A(\inv_in[1692] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1693] ));
 sky130_fd_sc_hd__inv_2 \inv[1693]/_0_  (.A(\inv_in[1693] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1694] ));
 sky130_fd_sc_hd__inv_2 \inv[1694]/_0_  (.A(\inv_in[1694] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1695] ));
 sky130_fd_sc_hd__inv_2 \inv[1695]/_0_  (.A(\inv_in[1695] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1696] ));
 sky130_fd_sc_hd__inv_2 \inv[1696]/_0_  (.A(\inv_in[1696] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1697] ));
 sky130_fd_sc_hd__inv_2 \inv[1697]/_0_  (.A(\inv_in[1697] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1698] ));
 sky130_fd_sc_hd__inv_2 \inv[1698]/_0_  (.A(\inv_in[1698] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1699] ));
 sky130_fd_sc_hd__inv_2 \inv[1699]/_0_  (.A(\inv_in[1699] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1700] ));
 sky130_fd_sc_hd__inv_2 \inv[169]/_0_  (.A(\inv_in[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[170] ));
 sky130_fd_sc_hd__inv_2 \inv[16]/_0_  (.A(\inv_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[17] ));
 sky130_fd_sc_hd__inv_2 \inv[1700]/_0_  (.A(\inv_in[1700] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1701] ));
 sky130_fd_sc_hd__inv_2 \inv[1701]/_0_  (.A(\inv_in[1701] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1702] ));
 sky130_fd_sc_hd__inv_2 \inv[1702]/_0_  (.A(\inv_in[1702] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1703] ));
 sky130_fd_sc_hd__inv_2 \inv[1703]/_0_  (.A(\inv_in[1703] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1704] ));
 sky130_fd_sc_hd__inv_2 \inv[1704]/_0_  (.A(\inv_in[1704] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1705] ));
 sky130_fd_sc_hd__inv_2 \inv[1705]/_0_  (.A(\inv_in[1705] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1706] ));
 sky130_fd_sc_hd__inv_2 \inv[1706]/_0_  (.A(\inv_in[1706] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1707] ));
 sky130_fd_sc_hd__inv_2 \inv[1707]/_0_  (.A(\inv_in[1707] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1708] ));
 sky130_fd_sc_hd__inv_2 \inv[1708]/_0_  (.A(\inv_in[1708] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1709] ));
 sky130_fd_sc_hd__inv_2 \inv[1709]/_0_  (.A(\inv_in[1709] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1710] ));
 sky130_fd_sc_hd__inv_2 \inv[170]/_0_  (.A(\inv_in[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[171] ));
 sky130_fd_sc_hd__inv_2 \inv[1710]/_0_  (.A(\inv_in[1710] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1711] ));
 sky130_fd_sc_hd__inv_2 \inv[1711]/_0_  (.A(\inv_in[1711] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1712] ));
 sky130_fd_sc_hd__inv_2 \inv[1712]/_0_  (.A(\inv_in[1712] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1713] ));
 sky130_fd_sc_hd__inv_2 \inv[1713]/_0_  (.A(\inv_in[1713] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1714] ));
 sky130_fd_sc_hd__inv_2 \inv[1714]/_0_  (.A(\inv_in[1714] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1715] ));
 sky130_fd_sc_hd__inv_2 \inv[1715]/_0_  (.A(\inv_in[1715] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1716] ));
 sky130_fd_sc_hd__inv_2 \inv[1716]/_0_  (.A(\inv_in[1716] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1717] ));
 sky130_fd_sc_hd__inv_2 \inv[1717]/_0_  (.A(\inv_in[1717] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1718] ));
 sky130_fd_sc_hd__inv_2 \inv[1718]/_0_  (.A(\inv_in[1718] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1719] ));
 sky130_fd_sc_hd__inv_2 \inv[1719]/_0_  (.A(\inv_in[1719] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1720] ));
 sky130_fd_sc_hd__inv_2 \inv[171]/_0_  (.A(\inv_in[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[172] ));
 sky130_fd_sc_hd__inv_2 \inv[1720]/_0_  (.A(\inv_in[1720] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1721] ));
 sky130_fd_sc_hd__inv_2 \inv[1721]/_0_  (.A(\inv_in[1721] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1722] ));
 sky130_fd_sc_hd__inv_2 \inv[1722]/_0_  (.A(\inv_in[1722] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1723] ));
 sky130_fd_sc_hd__inv_2 \inv[1723]/_0_  (.A(\inv_in[1723] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1724] ));
 sky130_fd_sc_hd__inv_2 \inv[1724]/_0_  (.A(\inv_in[1724] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1725] ));
 sky130_fd_sc_hd__inv_2 \inv[1725]/_0_  (.A(\inv_in[1725] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1726] ));
 sky130_fd_sc_hd__inv_2 \inv[1726]/_0_  (.A(\inv_in[1726] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1727] ));
 sky130_fd_sc_hd__inv_2 \inv[1727]/_0_  (.A(\inv_in[1727] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1728] ));
 sky130_fd_sc_hd__inv_2 \inv[1728]/_0_  (.A(\inv_in[1728] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1729] ));
 sky130_fd_sc_hd__inv_2 \inv[1729]/_0_  (.A(\inv_in[1729] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1730] ));
 sky130_fd_sc_hd__inv_2 \inv[172]/_0_  (.A(\inv_in[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[173] ));
 sky130_fd_sc_hd__inv_2 \inv[1730]/_0_  (.A(\inv_in[1730] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1731] ));
 sky130_fd_sc_hd__inv_2 \inv[1731]/_0_  (.A(\inv_in[1731] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1732] ));
 sky130_fd_sc_hd__inv_2 \inv[1732]/_0_  (.A(\inv_in[1732] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1733] ));
 sky130_fd_sc_hd__inv_2 \inv[1733]/_0_  (.A(\inv_in[1733] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1734] ));
 sky130_fd_sc_hd__inv_2 \inv[1734]/_0_  (.A(\inv_in[1734] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1735] ));
 sky130_fd_sc_hd__inv_2 \inv[1735]/_0_  (.A(\inv_in[1735] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1736] ));
 sky130_fd_sc_hd__inv_2 \inv[1736]/_0_  (.A(\inv_in[1736] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1737] ));
 sky130_fd_sc_hd__inv_2 \inv[1737]/_0_  (.A(\inv_in[1737] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1738] ));
 sky130_fd_sc_hd__inv_2 \inv[1738]/_0_  (.A(\inv_in[1738] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1739] ));
 sky130_fd_sc_hd__inv_2 \inv[1739]/_0_  (.A(\inv_in[1739] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1740] ));
 sky130_fd_sc_hd__inv_2 \inv[173]/_0_  (.A(\inv_in[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[174] ));
 sky130_fd_sc_hd__inv_2 \inv[1740]/_0_  (.A(\inv_in[1740] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1741] ));
 sky130_fd_sc_hd__inv_2 \inv[1741]/_0_  (.A(\inv_in[1741] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1742] ));
 sky130_fd_sc_hd__inv_2 \inv[1742]/_0_  (.A(\inv_in[1742] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1743] ));
 sky130_fd_sc_hd__inv_2 \inv[1743]/_0_  (.A(\inv_in[1743] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1744] ));
 sky130_fd_sc_hd__inv_2 \inv[1744]/_0_  (.A(\inv_in[1744] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1745] ));
 sky130_fd_sc_hd__inv_2 \inv[1745]/_0_  (.A(\inv_in[1745] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1746] ));
 sky130_fd_sc_hd__inv_2 \inv[1746]/_0_  (.A(\inv_in[1746] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1747] ));
 sky130_fd_sc_hd__inv_2 \inv[1747]/_0_  (.A(\inv_in[1747] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1748] ));
 sky130_fd_sc_hd__inv_2 \inv[1748]/_0_  (.A(\inv_in[1748] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1749] ));
 sky130_fd_sc_hd__inv_2 \inv[1749]/_0_  (.A(\inv_in[1749] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1750] ));
 sky130_fd_sc_hd__inv_2 \inv[174]/_0_  (.A(\inv_in[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[175] ));
 sky130_fd_sc_hd__inv_2 \inv[1750]/_0_  (.A(\inv_in[1750] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1751] ));
 sky130_fd_sc_hd__inv_2 \inv[1751]/_0_  (.A(\inv_in[1751] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1752] ));
 sky130_fd_sc_hd__inv_2 \inv[1752]/_0_  (.A(\inv_in[1752] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1753] ));
 sky130_fd_sc_hd__inv_2 \inv[1753]/_0_  (.A(\inv_in[1753] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1754] ));
 sky130_fd_sc_hd__inv_2 \inv[1754]/_0_  (.A(\inv_in[1754] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1755] ));
 sky130_fd_sc_hd__inv_2 \inv[1755]/_0_  (.A(\inv_in[1755] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1756] ));
 sky130_fd_sc_hd__inv_2 \inv[1756]/_0_  (.A(\inv_in[1756] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1757] ));
 sky130_fd_sc_hd__inv_2 \inv[1757]/_0_  (.A(\inv_in[1757] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1758] ));
 sky130_fd_sc_hd__inv_2 \inv[1758]/_0_  (.A(\inv_in[1758] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1759] ));
 sky130_fd_sc_hd__inv_2 \inv[1759]/_0_  (.A(\inv_in[1759] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1760] ));
 sky130_fd_sc_hd__inv_2 \inv[175]/_0_  (.A(\inv_in[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[176] ));
 sky130_fd_sc_hd__inv_2 \inv[1760]/_0_  (.A(\inv_in[1760] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1761] ));
 sky130_fd_sc_hd__inv_2 \inv[1761]/_0_  (.A(\inv_in[1761] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1762] ));
 sky130_fd_sc_hd__inv_2 \inv[1762]/_0_  (.A(\inv_in[1762] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1763] ));
 sky130_fd_sc_hd__inv_2 \inv[1763]/_0_  (.A(\inv_in[1763] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1764] ));
 sky130_fd_sc_hd__inv_2 \inv[1764]/_0_  (.A(\inv_in[1764] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1765] ));
 sky130_fd_sc_hd__inv_2 \inv[1765]/_0_  (.A(\inv_in[1765] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1766] ));
 sky130_fd_sc_hd__inv_2 \inv[1766]/_0_  (.A(\inv_in[1766] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1767] ));
 sky130_fd_sc_hd__inv_2 \inv[1767]/_0_  (.A(\inv_in[1767] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1768] ));
 sky130_fd_sc_hd__inv_2 \inv[1768]/_0_  (.A(\inv_in[1768] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1769] ));
 sky130_fd_sc_hd__inv_2 \inv[1769]/_0_  (.A(\inv_in[1769] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1770] ));
 sky130_fd_sc_hd__inv_2 \inv[176]/_0_  (.A(\inv_in[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[177] ));
 sky130_fd_sc_hd__inv_2 \inv[1770]/_0_  (.A(\inv_in[1770] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1771] ));
 sky130_fd_sc_hd__inv_2 \inv[1771]/_0_  (.A(\inv_in[1771] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1772] ));
 sky130_fd_sc_hd__inv_2 \inv[1772]/_0_  (.A(\inv_in[1772] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1773] ));
 sky130_fd_sc_hd__inv_2 \inv[1773]/_0_  (.A(\inv_in[1773] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1774] ));
 sky130_fd_sc_hd__inv_2 \inv[1774]/_0_  (.A(\inv_in[1774] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1775] ));
 sky130_fd_sc_hd__inv_2 \inv[1775]/_0_  (.A(\inv_in[1775] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1776] ));
 sky130_fd_sc_hd__inv_2 \inv[1776]/_0_  (.A(\inv_in[1776] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1777] ));
 sky130_fd_sc_hd__inv_2 \inv[1777]/_0_  (.A(\inv_in[1777] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1778] ));
 sky130_fd_sc_hd__inv_2 \inv[1778]/_0_  (.A(\inv_in[1778] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1779] ));
 sky130_fd_sc_hd__inv_2 \inv[1779]/_0_  (.A(\inv_in[1779] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1780] ));
 sky130_fd_sc_hd__inv_2 \inv[177]/_0_  (.A(\inv_in[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[178] ));
 sky130_fd_sc_hd__inv_2 \inv[1780]/_0_  (.A(\inv_in[1780] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1781] ));
 sky130_fd_sc_hd__inv_2 \inv[1781]/_0_  (.A(\inv_in[1781] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1782] ));
 sky130_fd_sc_hd__inv_2 \inv[1782]/_0_  (.A(\inv_in[1782] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1783] ));
 sky130_fd_sc_hd__inv_2 \inv[1783]/_0_  (.A(\inv_in[1783] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1784] ));
 sky130_fd_sc_hd__inv_2 \inv[1784]/_0_  (.A(\inv_in[1784] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1785] ));
 sky130_fd_sc_hd__inv_2 \inv[1785]/_0_  (.A(\inv_in[1785] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1786] ));
 sky130_fd_sc_hd__inv_2 \inv[1786]/_0_  (.A(\inv_in[1786] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1787] ));
 sky130_fd_sc_hd__inv_2 \inv[1787]/_0_  (.A(\inv_in[1787] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1788] ));
 sky130_fd_sc_hd__inv_2 \inv[1788]/_0_  (.A(\inv_in[1788] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1789] ));
 sky130_fd_sc_hd__inv_2 \inv[1789]/_0_  (.A(\inv_in[1789] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1790] ));
 sky130_fd_sc_hd__inv_2 \inv[178]/_0_  (.A(\inv_in[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[179] ));
 sky130_fd_sc_hd__inv_2 \inv[1790]/_0_  (.A(\inv_in[1790] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1791] ));
 sky130_fd_sc_hd__inv_2 \inv[1791]/_0_  (.A(\inv_in[1791] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1792] ));
 sky130_fd_sc_hd__inv_2 \inv[1792]/_0_  (.A(\inv_in[1792] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1793] ));
 sky130_fd_sc_hd__inv_2 \inv[1793]/_0_  (.A(\inv_in[1793] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1794] ));
 sky130_fd_sc_hd__inv_2 \inv[1794]/_0_  (.A(\inv_in[1794] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1795] ));
 sky130_fd_sc_hd__inv_2 \inv[1795]/_0_  (.A(\inv_in[1795] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1796] ));
 sky130_fd_sc_hd__inv_2 \inv[1796]/_0_  (.A(\inv_in[1796] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1797] ));
 sky130_fd_sc_hd__inv_2 \inv[1797]/_0_  (.A(\inv_in[1797] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1798] ));
 sky130_fd_sc_hd__inv_2 \inv[1798]/_0_  (.A(\inv_in[1798] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1799] ));
 sky130_fd_sc_hd__inv_2 \inv[1799]/_0_  (.A(\inv_in[1799] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1800] ));
 sky130_fd_sc_hd__inv_2 \inv[179]/_0_  (.A(\inv_in[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[180] ));
 sky130_fd_sc_hd__inv_2 \inv[17]/_0_  (.A(\inv_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[18] ));
 sky130_fd_sc_hd__inv_2 \inv[1800]/_0_  (.A(\inv_in[1800] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1801] ));
 sky130_fd_sc_hd__inv_2 \inv[1801]/_0_  (.A(\inv_in[1801] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1802] ));
 sky130_fd_sc_hd__inv_2 \inv[1802]/_0_  (.A(\inv_in[1802] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1803] ));
 sky130_fd_sc_hd__inv_2 \inv[1803]/_0_  (.A(\inv_in[1803] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1804] ));
 sky130_fd_sc_hd__inv_2 \inv[1804]/_0_  (.A(\inv_in[1804] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1805] ));
 sky130_fd_sc_hd__inv_2 \inv[1805]/_0_  (.A(\inv_in[1805] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1806] ));
 sky130_fd_sc_hd__inv_2 \inv[1806]/_0_  (.A(\inv_in[1806] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1807] ));
 sky130_fd_sc_hd__inv_2 \inv[1807]/_0_  (.A(\inv_in[1807] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1808] ));
 sky130_fd_sc_hd__inv_2 \inv[1808]/_0_  (.A(\inv_in[1808] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1809] ));
 sky130_fd_sc_hd__inv_2 \inv[1809]/_0_  (.A(\inv_in[1809] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1810] ));
 sky130_fd_sc_hd__inv_2 \inv[180]/_0_  (.A(\inv_in[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[181] ));
 sky130_fd_sc_hd__inv_2 \inv[1810]/_0_  (.A(\inv_in[1810] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1811] ));
 sky130_fd_sc_hd__inv_2 \inv[1811]/_0_  (.A(\inv_in[1811] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1812] ));
 sky130_fd_sc_hd__inv_2 \inv[1812]/_0_  (.A(\inv_in[1812] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1813] ));
 sky130_fd_sc_hd__inv_2 \inv[1813]/_0_  (.A(\inv_in[1813] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1814] ));
 sky130_fd_sc_hd__inv_2 \inv[1814]/_0_  (.A(\inv_in[1814] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1815] ));
 sky130_fd_sc_hd__inv_2 \inv[1815]/_0_  (.A(\inv_in[1815] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1816] ));
 sky130_fd_sc_hd__inv_2 \inv[1816]/_0_  (.A(\inv_in[1816] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1817] ));
 sky130_fd_sc_hd__inv_2 \inv[1817]/_0_  (.A(\inv_in[1817] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1818] ));
 sky130_fd_sc_hd__inv_2 \inv[1818]/_0_  (.A(\inv_in[1818] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1819] ));
 sky130_fd_sc_hd__inv_2 \inv[1819]/_0_  (.A(\inv_in[1819] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1820] ));
 sky130_fd_sc_hd__inv_2 \inv[181]/_0_  (.A(\inv_in[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[182] ));
 sky130_fd_sc_hd__inv_2 \inv[1820]/_0_  (.A(\inv_in[1820] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1821] ));
 sky130_fd_sc_hd__inv_2 \inv[1821]/_0_  (.A(\inv_in[1821] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1822] ));
 sky130_fd_sc_hd__inv_2 \inv[1822]/_0_  (.A(\inv_in[1822] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1823] ));
 sky130_fd_sc_hd__inv_2 \inv[1823]/_0_  (.A(\inv_in[1823] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1824] ));
 sky130_fd_sc_hd__inv_2 \inv[1824]/_0_  (.A(\inv_in[1824] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1825] ));
 sky130_fd_sc_hd__inv_2 \inv[1825]/_0_  (.A(\inv_in[1825] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1826] ));
 sky130_fd_sc_hd__inv_2 \inv[1826]/_0_  (.A(\inv_in[1826] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1827] ));
 sky130_fd_sc_hd__inv_2 \inv[1827]/_0_  (.A(\inv_in[1827] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1828] ));
 sky130_fd_sc_hd__inv_2 \inv[1828]/_0_  (.A(\inv_in[1828] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1829] ));
 sky130_fd_sc_hd__inv_2 \inv[1829]/_0_  (.A(\inv_in[1829] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1830] ));
 sky130_fd_sc_hd__inv_2 \inv[182]/_0_  (.A(\inv_in[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[183] ));
 sky130_fd_sc_hd__inv_2 \inv[1830]/_0_  (.A(\inv_in[1830] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1831] ));
 sky130_fd_sc_hd__inv_2 \inv[1831]/_0_  (.A(\inv_in[1831] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1832] ));
 sky130_fd_sc_hd__inv_2 \inv[1832]/_0_  (.A(\inv_in[1832] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1833] ));
 sky130_fd_sc_hd__inv_2 \inv[1833]/_0_  (.A(\inv_in[1833] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1834] ));
 sky130_fd_sc_hd__inv_2 \inv[1834]/_0_  (.A(\inv_in[1834] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1835] ));
 sky130_fd_sc_hd__inv_2 \inv[1835]/_0_  (.A(\inv_in[1835] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1836] ));
 sky130_fd_sc_hd__inv_2 \inv[1836]/_0_  (.A(\inv_in[1836] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1837] ));
 sky130_fd_sc_hd__inv_2 \inv[1837]/_0_  (.A(\inv_in[1837] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1838] ));
 sky130_fd_sc_hd__inv_2 \inv[1838]/_0_  (.A(\inv_in[1838] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1839] ));
 sky130_fd_sc_hd__inv_2 \inv[1839]/_0_  (.A(\inv_in[1839] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1840] ));
 sky130_fd_sc_hd__inv_2 \inv[183]/_0_  (.A(\inv_in[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[184] ));
 sky130_fd_sc_hd__inv_2 \inv[1840]/_0_  (.A(\inv_in[1840] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1841] ));
 sky130_fd_sc_hd__inv_2 \inv[1841]/_0_  (.A(\inv_in[1841] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1842] ));
 sky130_fd_sc_hd__inv_2 \inv[1842]/_0_  (.A(\inv_in[1842] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1843] ));
 sky130_fd_sc_hd__inv_2 \inv[1843]/_0_  (.A(\inv_in[1843] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1844] ));
 sky130_fd_sc_hd__inv_2 \inv[1844]/_0_  (.A(\inv_in[1844] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1845] ));
 sky130_fd_sc_hd__inv_2 \inv[1845]/_0_  (.A(\inv_in[1845] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1846] ));
 sky130_fd_sc_hd__inv_2 \inv[1846]/_0_  (.A(\inv_in[1846] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1847] ));
 sky130_fd_sc_hd__inv_2 \inv[1847]/_0_  (.A(\inv_in[1847] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1848] ));
 sky130_fd_sc_hd__inv_2 \inv[1848]/_0_  (.A(\inv_in[1848] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1849] ));
 sky130_fd_sc_hd__inv_2 \inv[1849]/_0_  (.A(\inv_in[1849] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1850] ));
 sky130_fd_sc_hd__inv_2 \inv[184]/_0_  (.A(\inv_in[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[185] ));
 sky130_fd_sc_hd__inv_2 \inv[1850]/_0_  (.A(\inv_in[1850] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1851] ));
 sky130_fd_sc_hd__inv_2 \inv[1851]/_0_  (.A(\inv_in[1851] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1852] ));
 sky130_fd_sc_hd__inv_2 \inv[1852]/_0_  (.A(\inv_in[1852] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1853] ));
 sky130_fd_sc_hd__inv_2 \inv[1853]/_0_  (.A(\inv_in[1853] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1854] ));
 sky130_fd_sc_hd__inv_2 \inv[1854]/_0_  (.A(\inv_in[1854] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1855] ));
 sky130_fd_sc_hd__inv_2 \inv[1855]/_0_  (.A(\inv_in[1855] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1856] ));
 sky130_fd_sc_hd__inv_2 \inv[1856]/_0_  (.A(\inv_in[1856] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1857] ));
 sky130_fd_sc_hd__inv_2 \inv[1857]/_0_  (.A(\inv_in[1857] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1858] ));
 sky130_fd_sc_hd__inv_2 \inv[1858]/_0_  (.A(\inv_in[1858] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1859] ));
 sky130_fd_sc_hd__inv_2 \inv[1859]/_0_  (.A(\inv_in[1859] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1860] ));
 sky130_fd_sc_hd__inv_2 \inv[185]/_0_  (.A(\inv_in[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[186] ));
 sky130_fd_sc_hd__inv_2 \inv[1860]/_0_  (.A(\inv_in[1860] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1861] ));
 sky130_fd_sc_hd__inv_2 \inv[1861]/_0_  (.A(\inv_in[1861] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1862] ));
 sky130_fd_sc_hd__inv_2 \inv[1862]/_0_  (.A(\inv_in[1862] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1863] ));
 sky130_fd_sc_hd__inv_2 \inv[1863]/_0_  (.A(\inv_in[1863] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1864] ));
 sky130_fd_sc_hd__inv_2 \inv[1864]/_0_  (.A(\inv_in[1864] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1865] ));
 sky130_fd_sc_hd__inv_2 \inv[1865]/_0_  (.A(\inv_in[1865] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1866] ));
 sky130_fd_sc_hd__inv_2 \inv[1866]/_0_  (.A(\inv_in[1866] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1867] ));
 sky130_fd_sc_hd__inv_2 \inv[1867]/_0_  (.A(\inv_in[1867] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1868] ));
 sky130_fd_sc_hd__inv_2 \inv[1868]/_0_  (.A(\inv_in[1868] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1869] ));
 sky130_fd_sc_hd__inv_2 \inv[1869]/_0_  (.A(\inv_in[1869] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1870] ));
 sky130_fd_sc_hd__inv_2 \inv[186]/_0_  (.A(\inv_in[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[187] ));
 sky130_fd_sc_hd__inv_2 \inv[1870]/_0_  (.A(\inv_in[1870] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1871] ));
 sky130_fd_sc_hd__inv_2 \inv[1871]/_0_  (.A(\inv_in[1871] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1872] ));
 sky130_fd_sc_hd__inv_2 \inv[1872]/_0_  (.A(\inv_in[1872] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1873] ));
 sky130_fd_sc_hd__inv_2 \inv[1873]/_0_  (.A(\inv_in[1873] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1874] ));
 sky130_fd_sc_hd__inv_2 \inv[1874]/_0_  (.A(\inv_in[1874] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1875] ));
 sky130_fd_sc_hd__inv_2 \inv[1875]/_0_  (.A(\inv_in[1875] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1876] ));
 sky130_fd_sc_hd__inv_2 \inv[1876]/_0_  (.A(\inv_in[1876] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1877] ));
 sky130_fd_sc_hd__inv_2 \inv[1877]/_0_  (.A(\inv_in[1877] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1878] ));
 sky130_fd_sc_hd__inv_2 \inv[1878]/_0_  (.A(\inv_in[1878] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1879] ));
 sky130_fd_sc_hd__inv_2 \inv[1879]/_0_  (.A(\inv_in[1879] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1880] ));
 sky130_fd_sc_hd__inv_2 \inv[187]/_0_  (.A(\inv_in[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[188] ));
 sky130_fd_sc_hd__inv_2 \inv[1880]/_0_  (.A(\inv_in[1880] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1881] ));
 sky130_fd_sc_hd__inv_2 \inv[1881]/_0_  (.A(\inv_in[1881] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1882] ));
 sky130_fd_sc_hd__inv_2 \inv[1882]/_0_  (.A(\inv_in[1882] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1883] ));
 sky130_fd_sc_hd__inv_2 \inv[1883]/_0_  (.A(\inv_in[1883] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1884] ));
 sky130_fd_sc_hd__inv_2 \inv[1884]/_0_  (.A(\inv_in[1884] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1885] ));
 sky130_fd_sc_hd__inv_2 \inv[1885]/_0_  (.A(\inv_in[1885] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1886] ));
 sky130_fd_sc_hd__inv_2 \inv[1886]/_0_  (.A(\inv_in[1886] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1887] ));
 sky130_fd_sc_hd__inv_2 \inv[1887]/_0_  (.A(\inv_in[1887] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1888] ));
 sky130_fd_sc_hd__inv_2 \inv[1888]/_0_  (.A(\inv_in[1888] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1889] ));
 sky130_fd_sc_hd__inv_2 \inv[1889]/_0_  (.A(\inv_in[1889] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1890] ));
 sky130_fd_sc_hd__inv_2 \inv[188]/_0_  (.A(\inv_in[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[189] ));
 sky130_fd_sc_hd__inv_2 \inv[1890]/_0_  (.A(\inv_in[1890] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1891] ));
 sky130_fd_sc_hd__inv_2 \inv[1891]/_0_  (.A(\inv_in[1891] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1892] ));
 sky130_fd_sc_hd__inv_2 \inv[1892]/_0_  (.A(\inv_in[1892] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1893] ));
 sky130_fd_sc_hd__inv_2 \inv[1893]/_0_  (.A(\inv_in[1893] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1894] ));
 sky130_fd_sc_hd__inv_2 \inv[1894]/_0_  (.A(\inv_in[1894] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1895] ));
 sky130_fd_sc_hd__inv_2 \inv[1895]/_0_  (.A(\inv_in[1895] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1896] ));
 sky130_fd_sc_hd__inv_2 \inv[1896]/_0_  (.A(\inv_in[1896] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1897] ));
 sky130_fd_sc_hd__inv_2 \inv[1897]/_0_  (.A(\inv_in[1897] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1898] ));
 sky130_fd_sc_hd__inv_2 \inv[1898]/_0_  (.A(\inv_in[1898] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1899] ));
 sky130_fd_sc_hd__inv_2 \inv[1899]/_0_  (.A(\inv_in[1899] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1900] ));
 sky130_fd_sc_hd__inv_2 \inv[189]/_0_  (.A(\inv_in[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[190] ));
 sky130_fd_sc_hd__inv_2 \inv[18]/_0_  (.A(\inv_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[19] ));
 sky130_fd_sc_hd__inv_2 \inv[1900]/_0_  (.A(\inv_in[1900] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1901] ));
 sky130_fd_sc_hd__inv_2 \inv[1901]/_0_  (.A(\inv_in[1901] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1902] ));
 sky130_fd_sc_hd__inv_2 \inv[1902]/_0_  (.A(\inv_in[1902] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1903] ));
 sky130_fd_sc_hd__inv_2 \inv[1903]/_0_  (.A(\inv_in[1903] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1904] ));
 sky130_fd_sc_hd__inv_2 \inv[1904]/_0_  (.A(\inv_in[1904] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1905] ));
 sky130_fd_sc_hd__inv_2 \inv[1905]/_0_  (.A(\inv_in[1905] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1906] ));
 sky130_fd_sc_hd__inv_2 \inv[1906]/_0_  (.A(\inv_in[1906] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1907] ));
 sky130_fd_sc_hd__inv_2 \inv[1907]/_0_  (.A(\inv_in[1907] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1908] ));
 sky130_fd_sc_hd__inv_2 \inv[1908]/_0_  (.A(\inv_in[1908] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1909] ));
 sky130_fd_sc_hd__inv_2 \inv[1909]/_0_  (.A(\inv_in[1909] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1910] ));
 sky130_fd_sc_hd__inv_2 \inv[190]/_0_  (.A(\inv_in[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[191] ));
 sky130_fd_sc_hd__inv_2 \inv[1910]/_0_  (.A(\inv_in[1910] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1911] ));
 sky130_fd_sc_hd__inv_2 \inv[1911]/_0_  (.A(\inv_in[1911] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1912] ));
 sky130_fd_sc_hd__inv_2 \inv[1912]/_0_  (.A(\inv_in[1912] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1913] ));
 sky130_fd_sc_hd__inv_2 \inv[1913]/_0_  (.A(\inv_in[1913] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1914] ));
 sky130_fd_sc_hd__inv_2 \inv[1914]/_0_  (.A(\inv_in[1914] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1915] ));
 sky130_fd_sc_hd__inv_2 \inv[1915]/_0_  (.A(\inv_in[1915] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1916] ));
 sky130_fd_sc_hd__inv_2 \inv[1916]/_0_  (.A(\inv_in[1916] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1917] ));
 sky130_fd_sc_hd__inv_2 \inv[1917]/_0_  (.A(\inv_in[1917] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1918] ));
 sky130_fd_sc_hd__inv_2 \inv[1918]/_0_  (.A(\inv_in[1918] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1919] ));
 sky130_fd_sc_hd__inv_2 \inv[1919]/_0_  (.A(\inv_in[1919] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1920] ));
 sky130_fd_sc_hd__inv_2 \inv[191]/_0_  (.A(\inv_in[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[192] ));
 sky130_fd_sc_hd__inv_2 \inv[1920]/_0_  (.A(\inv_in[1920] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1921] ));
 sky130_fd_sc_hd__inv_2 \inv[1921]/_0_  (.A(\inv_in[1921] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1922] ));
 sky130_fd_sc_hd__inv_2 \inv[1922]/_0_  (.A(\inv_in[1922] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1923] ));
 sky130_fd_sc_hd__inv_2 \inv[1923]/_0_  (.A(\inv_in[1923] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1924] ));
 sky130_fd_sc_hd__inv_2 \inv[1924]/_0_  (.A(\inv_in[1924] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1925] ));
 sky130_fd_sc_hd__inv_2 \inv[1925]/_0_  (.A(\inv_in[1925] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1926] ));
 sky130_fd_sc_hd__inv_2 \inv[1926]/_0_  (.A(\inv_in[1926] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1927] ));
 sky130_fd_sc_hd__inv_2 \inv[1927]/_0_  (.A(\inv_in[1927] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1928] ));
 sky130_fd_sc_hd__inv_2 \inv[1928]/_0_  (.A(\inv_in[1928] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1929] ));
 sky130_fd_sc_hd__inv_2 \inv[1929]/_0_  (.A(\inv_in[1929] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1930] ));
 sky130_fd_sc_hd__inv_2 \inv[192]/_0_  (.A(\inv_in[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[193] ));
 sky130_fd_sc_hd__inv_2 \inv[1930]/_0_  (.A(\inv_in[1930] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1931] ));
 sky130_fd_sc_hd__inv_2 \inv[1931]/_0_  (.A(\inv_in[1931] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1932] ));
 sky130_fd_sc_hd__inv_2 \inv[1932]/_0_  (.A(\inv_in[1932] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1933] ));
 sky130_fd_sc_hd__inv_2 \inv[1933]/_0_  (.A(\inv_in[1933] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1934] ));
 sky130_fd_sc_hd__inv_2 \inv[1934]/_0_  (.A(\inv_in[1934] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1935] ));
 sky130_fd_sc_hd__inv_2 \inv[1935]/_0_  (.A(\inv_in[1935] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1936] ));
 sky130_fd_sc_hd__inv_2 \inv[1936]/_0_  (.A(\inv_in[1936] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1937] ));
 sky130_fd_sc_hd__inv_2 \inv[1937]/_0_  (.A(\inv_in[1937] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1938] ));
 sky130_fd_sc_hd__inv_2 \inv[1938]/_0_  (.A(\inv_in[1938] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1939] ));
 sky130_fd_sc_hd__inv_2 \inv[1939]/_0_  (.A(\inv_in[1939] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1940] ));
 sky130_fd_sc_hd__inv_2 \inv[193]/_0_  (.A(\inv_in[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[194] ));
 sky130_fd_sc_hd__inv_2 \inv[1940]/_0_  (.A(\inv_in[1940] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1941] ));
 sky130_fd_sc_hd__inv_2 \inv[1941]/_0_  (.A(\inv_in[1941] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1942] ));
 sky130_fd_sc_hd__inv_2 \inv[1942]/_0_  (.A(\inv_in[1942] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1943] ));
 sky130_fd_sc_hd__inv_2 \inv[1943]/_0_  (.A(\inv_in[1943] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1944] ));
 sky130_fd_sc_hd__inv_2 \inv[1944]/_0_  (.A(\inv_in[1944] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1945] ));
 sky130_fd_sc_hd__inv_2 \inv[1945]/_0_  (.A(\inv_in[1945] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1946] ));
 sky130_fd_sc_hd__inv_2 \inv[1946]/_0_  (.A(\inv_in[1946] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1947] ));
 sky130_fd_sc_hd__inv_2 \inv[1947]/_0_  (.A(\inv_in[1947] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1948] ));
 sky130_fd_sc_hd__inv_2 \inv[1948]/_0_  (.A(\inv_in[1948] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1949] ));
 sky130_fd_sc_hd__inv_2 \inv[1949]/_0_  (.A(\inv_in[1949] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1950] ));
 sky130_fd_sc_hd__inv_2 \inv[194]/_0_  (.A(\inv_in[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[195] ));
 sky130_fd_sc_hd__inv_2 \inv[1950]/_0_  (.A(\inv_in[1950] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1951] ));
 sky130_fd_sc_hd__inv_2 \inv[1951]/_0_  (.A(\inv_in[1951] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1952] ));
 sky130_fd_sc_hd__inv_2 \inv[1952]/_0_  (.A(\inv_in[1952] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1953] ));
 sky130_fd_sc_hd__inv_2 \inv[1953]/_0_  (.A(\inv_in[1953] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1954] ));
 sky130_fd_sc_hd__inv_2 \inv[1954]/_0_  (.A(\inv_in[1954] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1955] ));
 sky130_fd_sc_hd__inv_2 \inv[1955]/_0_  (.A(\inv_in[1955] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1956] ));
 sky130_fd_sc_hd__inv_2 \inv[1956]/_0_  (.A(\inv_in[1956] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1957] ));
 sky130_fd_sc_hd__inv_2 \inv[1957]/_0_  (.A(\inv_in[1957] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1958] ));
 sky130_fd_sc_hd__inv_2 \inv[1958]/_0_  (.A(\inv_in[1958] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1959] ));
 sky130_fd_sc_hd__inv_2 \inv[1959]/_0_  (.A(\inv_in[1959] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1960] ));
 sky130_fd_sc_hd__inv_2 \inv[195]/_0_  (.A(\inv_in[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[196] ));
 sky130_fd_sc_hd__inv_2 \inv[1960]/_0_  (.A(\inv_in[1960] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1961] ));
 sky130_fd_sc_hd__inv_2 \inv[1961]/_0_  (.A(\inv_in[1961] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1962] ));
 sky130_fd_sc_hd__inv_2 \inv[1962]/_0_  (.A(\inv_in[1962] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1963] ));
 sky130_fd_sc_hd__inv_2 \inv[1963]/_0_  (.A(\inv_in[1963] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1964] ));
 sky130_fd_sc_hd__inv_2 \inv[1964]/_0_  (.A(\inv_in[1964] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1965] ));
 sky130_fd_sc_hd__inv_2 \inv[1965]/_0_  (.A(\inv_in[1965] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1966] ));
 sky130_fd_sc_hd__inv_2 \inv[1966]/_0_  (.A(\inv_in[1966] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1967] ));
 sky130_fd_sc_hd__inv_2 \inv[1967]/_0_  (.A(\inv_in[1967] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1968] ));
 sky130_fd_sc_hd__inv_2 \inv[1968]/_0_  (.A(\inv_in[1968] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1969] ));
 sky130_fd_sc_hd__inv_2 \inv[1969]/_0_  (.A(\inv_in[1969] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1970] ));
 sky130_fd_sc_hd__inv_2 \inv[196]/_0_  (.A(\inv_in[196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[197] ));
 sky130_fd_sc_hd__inv_2 \inv[1970]/_0_  (.A(\inv_in[1970] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1971] ));
 sky130_fd_sc_hd__inv_2 \inv[1971]/_0_  (.A(\inv_in[1971] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1972] ));
 sky130_fd_sc_hd__inv_2 \inv[1972]/_0_  (.A(\inv_in[1972] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1973] ));
 sky130_fd_sc_hd__inv_2 \inv[1973]/_0_  (.A(\inv_in[1973] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1974] ));
 sky130_fd_sc_hd__inv_2 \inv[1974]/_0_  (.A(\inv_in[1974] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1975] ));
 sky130_fd_sc_hd__inv_2 \inv[1975]/_0_  (.A(\inv_in[1975] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1976] ));
 sky130_fd_sc_hd__inv_2 \inv[1976]/_0_  (.A(\inv_in[1976] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1977] ));
 sky130_fd_sc_hd__inv_2 \inv[1977]/_0_  (.A(\inv_in[1977] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1978] ));
 sky130_fd_sc_hd__inv_2 \inv[1978]/_0_  (.A(\inv_in[1978] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1979] ));
 sky130_fd_sc_hd__inv_2 \inv[1979]/_0_  (.A(\inv_in[1979] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1980] ));
 sky130_fd_sc_hd__inv_2 \inv[197]/_0_  (.A(\inv_in[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[198] ));
 sky130_fd_sc_hd__inv_2 \inv[1980]/_0_  (.A(\inv_in[1980] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1981] ));
 sky130_fd_sc_hd__inv_2 \inv[1981]/_0_  (.A(\inv_in[1981] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1982] ));
 sky130_fd_sc_hd__inv_2 \inv[1982]/_0_  (.A(\inv_in[1982] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1983] ));
 sky130_fd_sc_hd__inv_2 \inv[1983]/_0_  (.A(\inv_in[1983] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1984] ));
 sky130_fd_sc_hd__inv_2 \inv[1984]/_0_  (.A(\inv_in[1984] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1985] ));
 sky130_fd_sc_hd__inv_2 \inv[1985]/_0_  (.A(\inv_in[1985] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1986] ));
 sky130_fd_sc_hd__inv_2 \inv[1986]/_0_  (.A(\inv_in[1986] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1987] ));
 sky130_fd_sc_hd__inv_2 \inv[1987]/_0_  (.A(\inv_in[1987] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1988] ));
 sky130_fd_sc_hd__inv_2 \inv[1988]/_0_  (.A(\inv_in[1988] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1989] ));
 sky130_fd_sc_hd__inv_2 \inv[1989]/_0_  (.A(\inv_in[1989] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1990] ));
 sky130_fd_sc_hd__inv_2 \inv[198]/_0_  (.A(\inv_in[198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[199] ));
 sky130_fd_sc_hd__inv_2 \inv[1990]/_0_  (.A(\inv_in[1990] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1991] ));
 sky130_fd_sc_hd__inv_2 \inv[1991]/_0_  (.A(\inv_in[1991] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1992] ));
 sky130_fd_sc_hd__inv_2 \inv[1992]/_0_  (.A(\inv_in[1992] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1993] ));
 sky130_fd_sc_hd__inv_2 \inv[1993]/_0_  (.A(\inv_in[1993] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1994] ));
 sky130_fd_sc_hd__inv_2 \inv[1994]/_0_  (.A(\inv_in[1994] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1995] ));
 sky130_fd_sc_hd__inv_2 \inv[1995]/_0_  (.A(\inv_in[1995] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1996] ));
 sky130_fd_sc_hd__inv_2 \inv[1996]/_0_  (.A(\inv_in[1996] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1997] ));
 sky130_fd_sc_hd__inv_2 \inv[1997]/_0_  (.A(\inv_in[1997] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1998] ));
 sky130_fd_sc_hd__inv_2 \inv[1998]/_0_  (.A(\inv_in[1998] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1999] ));
 sky130_fd_sc_hd__inv_2 \inv[1999]/_0_  (.A(\inv_in[1999] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2000] ));
 sky130_fd_sc_hd__inv_2 \inv[199]/_0_  (.A(\inv_in[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[200] ));
 sky130_fd_sc_hd__inv_2 \inv[19]/_0_  (.A(\inv_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[20] ));
 sky130_fd_sc_hd__inv_2 \inv[1]/_0_  (.A(\inv_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2] ));
 sky130_fd_sc_hd__inv_2 \inv[2000]/_0_  (.A(\inv_in[2000] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2001] ));
 sky130_fd_sc_hd__inv_2 \inv[2001]/_0_  (.A(\inv_in[2001] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2002] ));
 sky130_fd_sc_hd__inv_2 \inv[2002]/_0_  (.A(\inv_in[2002] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2003] ));
 sky130_fd_sc_hd__inv_2 \inv[2003]/_0_  (.A(\inv_in[2003] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2004] ));
 sky130_fd_sc_hd__inv_2 \inv[2004]/_0_  (.A(\inv_in[2004] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2005] ));
 sky130_fd_sc_hd__inv_2 \inv[2005]/_0_  (.A(\inv_in[2005] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2006] ));
 sky130_fd_sc_hd__inv_2 \inv[2006]/_0_  (.A(\inv_in[2006] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2007] ));
 sky130_fd_sc_hd__inv_2 \inv[2007]/_0_  (.A(\inv_in[2007] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2008] ));
 sky130_fd_sc_hd__inv_2 \inv[2008]/_0_  (.A(\inv_in[2008] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2009] ));
 sky130_fd_sc_hd__inv_2 \inv[2009]/_0_  (.A(\inv_in[2009] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2010] ));
 sky130_fd_sc_hd__inv_2 \inv[200]/_0_  (.A(\inv_in[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[201] ));
 sky130_fd_sc_hd__inv_2 \inv[2010]/_0_  (.A(\inv_in[2010] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2011] ));
 sky130_fd_sc_hd__inv_2 \inv[2011]/_0_  (.A(\inv_in[2011] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2012] ));
 sky130_fd_sc_hd__inv_2 \inv[2012]/_0_  (.A(\inv_in[2012] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2013] ));
 sky130_fd_sc_hd__inv_2 \inv[2013]/_0_  (.A(\inv_in[2013] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2014] ));
 sky130_fd_sc_hd__inv_2 \inv[2014]/_0_  (.A(\inv_in[2014] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2015] ));
 sky130_fd_sc_hd__inv_2 \inv[2015]/_0_  (.A(\inv_in[2015] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2016] ));
 sky130_fd_sc_hd__inv_2 \inv[2016]/_0_  (.A(\inv_in[2016] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2017] ));
 sky130_fd_sc_hd__inv_2 \inv[2017]/_0_  (.A(\inv_in[2017] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2018] ));
 sky130_fd_sc_hd__inv_2 \inv[2018]/_0_  (.A(\inv_in[2018] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2019] ));
 sky130_fd_sc_hd__inv_2 \inv[2019]/_0_  (.A(\inv_in[2019] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2020] ));
 sky130_fd_sc_hd__inv_2 \inv[201]/_0_  (.A(\inv_in[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[202] ));
 sky130_fd_sc_hd__inv_2 \inv[2020]/_0_  (.A(\inv_in[2020] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2021] ));
 sky130_fd_sc_hd__inv_2 \inv[2021]/_0_  (.A(\inv_in[2021] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2022] ));
 sky130_fd_sc_hd__inv_2 \inv[2022]/_0_  (.A(\inv_in[2022] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2023] ));
 sky130_fd_sc_hd__inv_2 \inv[2023]/_0_  (.A(\inv_in[2023] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2024] ));
 sky130_fd_sc_hd__inv_2 \inv[2024]/_0_  (.A(\inv_in[2024] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2025] ));
 sky130_fd_sc_hd__inv_2 \inv[2025]/_0_  (.A(\inv_in[2025] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2026] ));
 sky130_fd_sc_hd__inv_2 \inv[2026]/_0_  (.A(\inv_in[2026] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2027] ));
 sky130_fd_sc_hd__inv_2 \inv[2027]/_0_  (.A(\inv_in[2027] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2028] ));
 sky130_fd_sc_hd__inv_2 \inv[2028]/_0_  (.A(\inv_in[2028] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2029] ));
 sky130_fd_sc_hd__inv_2 \inv[2029]/_0_  (.A(\inv_in[2029] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2030] ));
 sky130_fd_sc_hd__inv_2 \inv[202]/_0_  (.A(\inv_in[202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[203] ));
 sky130_fd_sc_hd__inv_2 \inv[2030]/_0_  (.A(\inv_in[2030] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2031] ));
 sky130_fd_sc_hd__inv_2 \inv[2031]/_0_  (.A(\inv_in[2031] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2032] ));
 sky130_fd_sc_hd__inv_2 \inv[2032]/_0_  (.A(\inv_in[2032] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2033] ));
 sky130_fd_sc_hd__inv_2 \inv[2033]/_0_  (.A(\inv_in[2033] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2034] ));
 sky130_fd_sc_hd__inv_2 \inv[2034]/_0_  (.A(\inv_in[2034] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2035] ));
 sky130_fd_sc_hd__inv_2 \inv[2035]/_0_  (.A(\inv_in[2035] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2036] ));
 sky130_fd_sc_hd__inv_2 \inv[2036]/_0_  (.A(\inv_in[2036] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2037] ));
 sky130_fd_sc_hd__inv_2 \inv[2037]/_0_  (.A(\inv_in[2037] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2038] ));
 sky130_fd_sc_hd__inv_2 \inv[2038]/_0_  (.A(\inv_in[2038] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2039] ));
 sky130_fd_sc_hd__inv_2 \inv[2039]/_0_  (.A(\inv_in[2039] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2040] ));
 sky130_fd_sc_hd__inv_2 \inv[203]/_0_  (.A(\inv_in[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[204] ));
 sky130_fd_sc_hd__inv_2 \inv[2040]/_0_  (.A(\inv_in[2040] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2041] ));
 sky130_fd_sc_hd__inv_2 \inv[2041]/_0_  (.A(\inv_in[2041] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2042] ));
 sky130_fd_sc_hd__inv_2 \inv[2042]/_0_  (.A(\inv_in[2042] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2043] ));
 sky130_fd_sc_hd__inv_2 \inv[2043]/_0_  (.A(\inv_in[2043] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2044] ));
 sky130_fd_sc_hd__inv_2 \inv[2044]/_0_  (.A(\inv_in[2044] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2045] ));
 sky130_fd_sc_hd__inv_2 \inv[2045]/_0_  (.A(\inv_in[2045] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2046] ));
 sky130_fd_sc_hd__inv_2 \inv[2046]/_0_  (.A(\inv_in[2046] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2047] ));
 sky130_fd_sc_hd__inv_2 \inv[2047]/_0_  (.A(\inv_in[2047] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2048] ));
 sky130_fd_sc_hd__inv_2 \inv[2048]/_0_  (.A(\inv_in[2048] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2049] ));
 sky130_fd_sc_hd__inv_2 \inv[2049]/_0_  (.A(\inv_in[2049] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2050] ));
 sky130_fd_sc_hd__inv_2 \inv[204]/_0_  (.A(\inv_in[204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[205] ));
 sky130_fd_sc_hd__inv_2 \inv[2050]/_0_  (.A(\inv_in[2050] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2051] ));
 sky130_fd_sc_hd__inv_2 \inv[2051]/_0_  (.A(\inv_in[2051] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2052] ));
 sky130_fd_sc_hd__inv_2 \inv[2052]/_0_  (.A(\inv_in[2052] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2053] ));
 sky130_fd_sc_hd__inv_2 \inv[2053]/_0_  (.A(\inv_in[2053] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2054] ));
 sky130_fd_sc_hd__inv_2 \inv[2054]/_0_  (.A(\inv_in[2054] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2055] ));
 sky130_fd_sc_hd__inv_2 \inv[2055]/_0_  (.A(\inv_in[2055] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2056] ));
 sky130_fd_sc_hd__inv_2 \inv[2056]/_0_  (.A(\inv_in[2056] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2057] ));
 sky130_fd_sc_hd__inv_2 \inv[2057]/_0_  (.A(\inv_in[2057] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2058] ));
 sky130_fd_sc_hd__inv_2 \inv[2058]/_0_  (.A(\inv_in[2058] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2059] ));
 sky130_fd_sc_hd__inv_2 \inv[2059]/_0_  (.A(\inv_in[2059] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2060] ));
 sky130_fd_sc_hd__inv_2 \inv[205]/_0_  (.A(\inv_in[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[206] ));
 sky130_fd_sc_hd__inv_2 \inv[2060]/_0_  (.A(\inv_in[2060] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2061] ));
 sky130_fd_sc_hd__inv_2 \inv[2061]/_0_  (.A(\inv_in[2061] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2062] ));
 sky130_fd_sc_hd__inv_2 \inv[2062]/_0_  (.A(\inv_in[2062] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2063] ));
 sky130_fd_sc_hd__inv_2 \inv[2063]/_0_  (.A(\inv_in[2063] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2064] ));
 sky130_fd_sc_hd__inv_2 \inv[2064]/_0_  (.A(\inv_in[2064] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2065] ));
 sky130_fd_sc_hd__inv_2 \inv[2065]/_0_  (.A(\inv_in[2065] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2066] ));
 sky130_fd_sc_hd__inv_2 \inv[2066]/_0_  (.A(\inv_in[2066] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2067] ));
 sky130_fd_sc_hd__inv_2 \inv[2067]/_0_  (.A(\inv_in[2067] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2068] ));
 sky130_fd_sc_hd__inv_2 \inv[2068]/_0_  (.A(\inv_in[2068] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2069] ));
 sky130_fd_sc_hd__inv_2 \inv[2069]/_0_  (.A(\inv_in[2069] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2070] ));
 sky130_fd_sc_hd__inv_2 \inv[206]/_0_  (.A(\inv_in[206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[207] ));
 sky130_fd_sc_hd__inv_2 \inv[2070]/_0_  (.A(\inv_in[2070] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2071] ));
 sky130_fd_sc_hd__inv_2 \inv[2071]/_0_  (.A(\inv_in[2071] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2072] ));
 sky130_fd_sc_hd__inv_2 \inv[2072]/_0_  (.A(\inv_in[2072] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2073] ));
 sky130_fd_sc_hd__inv_2 \inv[2073]/_0_  (.A(\inv_in[2073] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2074] ));
 sky130_fd_sc_hd__inv_2 \inv[2074]/_0_  (.A(\inv_in[2074] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2075] ));
 sky130_fd_sc_hd__inv_2 \inv[2075]/_0_  (.A(\inv_in[2075] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2076] ));
 sky130_fd_sc_hd__inv_2 \inv[2076]/_0_  (.A(\inv_in[2076] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2077] ));
 sky130_fd_sc_hd__inv_2 \inv[2077]/_0_  (.A(\inv_in[2077] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2078] ));
 sky130_fd_sc_hd__inv_2 \inv[2078]/_0_  (.A(\inv_in[2078] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2079] ));
 sky130_fd_sc_hd__inv_2 \inv[2079]/_0_  (.A(\inv_in[2079] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2080] ));
 sky130_fd_sc_hd__inv_2 \inv[207]/_0_  (.A(\inv_in[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[208] ));
 sky130_fd_sc_hd__inv_2 \inv[2080]/_0_  (.A(\inv_in[2080] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2081] ));
 sky130_fd_sc_hd__inv_2 \inv[2081]/_0_  (.A(\inv_in[2081] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2082] ));
 sky130_fd_sc_hd__inv_2 \inv[2082]/_0_  (.A(\inv_in[2082] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2083] ));
 sky130_fd_sc_hd__inv_2 \inv[2083]/_0_  (.A(\inv_in[2083] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2084] ));
 sky130_fd_sc_hd__inv_2 \inv[2084]/_0_  (.A(\inv_in[2084] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2085] ));
 sky130_fd_sc_hd__inv_2 \inv[2085]/_0_  (.A(\inv_in[2085] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2086] ));
 sky130_fd_sc_hd__inv_2 \inv[2086]/_0_  (.A(\inv_in[2086] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2087] ));
 sky130_fd_sc_hd__inv_2 \inv[2087]/_0_  (.A(\inv_in[2087] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2088] ));
 sky130_fd_sc_hd__inv_2 \inv[2088]/_0_  (.A(\inv_in[2088] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2089] ));
 sky130_fd_sc_hd__inv_2 \inv[2089]/_0_  (.A(\inv_in[2089] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2090] ));
 sky130_fd_sc_hd__inv_2 \inv[208]/_0_  (.A(\inv_in[208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[209] ));
 sky130_fd_sc_hd__inv_2 \inv[2090]/_0_  (.A(\inv_in[2090] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2091] ));
 sky130_fd_sc_hd__inv_2 \inv[2091]/_0_  (.A(\inv_in[2091] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2092] ));
 sky130_fd_sc_hd__inv_2 \inv[2092]/_0_  (.A(\inv_in[2092] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2093] ));
 sky130_fd_sc_hd__inv_2 \inv[2093]/_0_  (.A(\inv_in[2093] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2094] ));
 sky130_fd_sc_hd__inv_2 \inv[2094]/_0_  (.A(\inv_in[2094] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2095] ));
 sky130_fd_sc_hd__inv_2 \inv[2095]/_0_  (.A(\inv_in[2095] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2096] ));
 sky130_fd_sc_hd__inv_2 \inv[2096]/_0_  (.A(\inv_in[2096] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2097] ));
 sky130_fd_sc_hd__inv_2 \inv[2097]/_0_  (.A(\inv_in[2097] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2098] ));
 sky130_fd_sc_hd__inv_2 \inv[2098]/_0_  (.A(\inv_in[2098] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2099] ));
 sky130_fd_sc_hd__inv_2 \inv[2099]/_0_  (.A(\inv_in[2099] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2100] ));
 sky130_fd_sc_hd__inv_2 \inv[209]/_0_  (.A(\inv_in[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[210] ));
 sky130_fd_sc_hd__inv_2 \inv[20]/_0_  (.A(\inv_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[21] ));
 sky130_fd_sc_hd__inv_2 \inv[2100]/_0_  (.A(\inv_in[2100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2101] ));
 sky130_fd_sc_hd__inv_2 \inv[2101]/_0_  (.A(\inv_in[2101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2102] ));
 sky130_fd_sc_hd__inv_2 \inv[2102]/_0_  (.A(\inv_in[2102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2103] ));
 sky130_fd_sc_hd__inv_2 \inv[2103]/_0_  (.A(\inv_in[2103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2104] ));
 sky130_fd_sc_hd__inv_2 \inv[2104]/_0_  (.A(\inv_in[2104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2105] ));
 sky130_fd_sc_hd__inv_2 \inv[2105]/_0_  (.A(\inv_in[2105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2106] ));
 sky130_fd_sc_hd__inv_2 \inv[2106]/_0_  (.A(\inv_in[2106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2107] ));
 sky130_fd_sc_hd__inv_2 \inv[2107]/_0_  (.A(\inv_in[2107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2108] ));
 sky130_fd_sc_hd__inv_2 \inv[2108]/_0_  (.A(\inv_in[2108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2109] ));
 sky130_fd_sc_hd__inv_2 \inv[2109]/_0_  (.A(\inv_in[2109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2110] ));
 sky130_fd_sc_hd__inv_2 \inv[210]/_0_  (.A(\inv_in[210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[211] ));
 sky130_fd_sc_hd__inv_2 \inv[2110]/_0_  (.A(\inv_in[2110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2111] ));
 sky130_fd_sc_hd__inv_2 \inv[2111]/_0_  (.A(\inv_in[2111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2112] ));
 sky130_fd_sc_hd__inv_2 \inv[2112]/_0_  (.A(\inv_in[2112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2113] ));
 sky130_fd_sc_hd__inv_2 \inv[2113]/_0_  (.A(\inv_in[2113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2114] ));
 sky130_fd_sc_hd__inv_2 \inv[2114]/_0_  (.A(\inv_in[2114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2115] ));
 sky130_fd_sc_hd__inv_2 \inv[2115]/_0_  (.A(\inv_in[2115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2116] ));
 sky130_fd_sc_hd__inv_2 \inv[2116]/_0_  (.A(\inv_in[2116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2117] ));
 sky130_fd_sc_hd__inv_2 \inv[2117]/_0_  (.A(\inv_in[2117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2118] ));
 sky130_fd_sc_hd__inv_2 \inv[2118]/_0_  (.A(\inv_in[2118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2119] ));
 sky130_fd_sc_hd__inv_2 \inv[2119]/_0_  (.A(\inv_in[2119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2120] ));
 sky130_fd_sc_hd__inv_2 \inv[211]/_0_  (.A(\inv_in[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[212] ));
 sky130_fd_sc_hd__inv_2 \inv[2120]/_0_  (.A(\inv_in[2120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2121] ));
 sky130_fd_sc_hd__inv_2 \inv[2121]/_0_  (.A(\inv_in[2121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2122] ));
 sky130_fd_sc_hd__inv_2 \inv[2122]/_0_  (.A(\inv_in[2122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2123] ));
 sky130_fd_sc_hd__inv_2 \inv[2123]/_0_  (.A(\inv_in[2123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2124] ));
 sky130_fd_sc_hd__inv_2 \inv[2124]/_0_  (.A(\inv_in[2124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2125] ));
 sky130_fd_sc_hd__inv_2 \inv[2125]/_0_  (.A(\inv_in[2125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2126] ));
 sky130_fd_sc_hd__inv_2 \inv[2126]/_0_  (.A(\inv_in[2126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2127] ));
 sky130_fd_sc_hd__inv_2 \inv[2127]/_0_  (.A(\inv_in[2127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2128] ));
 sky130_fd_sc_hd__inv_2 \inv[2128]/_0_  (.A(\inv_in[2128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2129] ));
 sky130_fd_sc_hd__inv_2 \inv[2129]/_0_  (.A(\inv_in[2129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2130] ));
 sky130_fd_sc_hd__inv_2 \inv[212]/_0_  (.A(\inv_in[212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[213] ));
 sky130_fd_sc_hd__inv_2 \inv[2130]/_0_  (.A(\inv_in[2130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2131] ));
 sky130_fd_sc_hd__inv_2 \inv[2131]/_0_  (.A(\inv_in[2131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2132] ));
 sky130_fd_sc_hd__inv_2 \inv[2132]/_0_  (.A(\inv_in[2132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2133] ));
 sky130_fd_sc_hd__inv_2 \inv[2133]/_0_  (.A(\inv_in[2133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2134] ));
 sky130_fd_sc_hd__inv_2 \inv[2134]/_0_  (.A(\inv_in[2134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2135] ));
 sky130_fd_sc_hd__inv_2 \inv[2135]/_0_  (.A(\inv_in[2135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2136] ));
 sky130_fd_sc_hd__inv_2 \inv[2136]/_0_  (.A(\inv_in[2136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2137] ));
 sky130_fd_sc_hd__inv_2 \inv[2137]/_0_  (.A(\inv_in[2137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2138] ));
 sky130_fd_sc_hd__inv_2 \inv[2138]/_0_  (.A(\inv_in[2138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2139] ));
 sky130_fd_sc_hd__inv_2 \inv[2139]/_0_  (.A(\inv_in[2139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2140] ));
 sky130_fd_sc_hd__inv_2 \inv[213]/_0_  (.A(\inv_in[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[214] ));
 sky130_fd_sc_hd__inv_2 \inv[2140]/_0_  (.A(\inv_in[2140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2141] ));
 sky130_fd_sc_hd__inv_2 \inv[2141]/_0_  (.A(\inv_in[2141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2142] ));
 sky130_fd_sc_hd__inv_2 \inv[2142]/_0_  (.A(\inv_in[2142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2143] ));
 sky130_fd_sc_hd__inv_2 \inv[2143]/_0_  (.A(\inv_in[2143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2144] ));
 sky130_fd_sc_hd__inv_2 \inv[2144]/_0_  (.A(\inv_in[2144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2145] ));
 sky130_fd_sc_hd__inv_2 \inv[2145]/_0_  (.A(\inv_in[2145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2146] ));
 sky130_fd_sc_hd__inv_2 \inv[2146]/_0_  (.A(\inv_in[2146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2147] ));
 sky130_fd_sc_hd__inv_2 \inv[2147]/_0_  (.A(\inv_in[2147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2148] ));
 sky130_fd_sc_hd__inv_2 \inv[2148]/_0_  (.A(\inv_in[2148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2149] ));
 sky130_fd_sc_hd__inv_2 \inv[2149]/_0_  (.A(\inv_in[2149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2150] ));
 sky130_fd_sc_hd__inv_2 \inv[214]/_0_  (.A(\inv_in[214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[215] ));
 sky130_fd_sc_hd__inv_2 \inv[2150]/_0_  (.A(\inv_in[2150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2151] ));
 sky130_fd_sc_hd__inv_2 \inv[2151]/_0_  (.A(\inv_in[2151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2152] ));
 sky130_fd_sc_hd__inv_2 \inv[2152]/_0_  (.A(\inv_in[2152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2153] ));
 sky130_fd_sc_hd__inv_2 \inv[2153]/_0_  (.A(\inv_in[2153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2154] ));
 sky130_fd_sc_hd__inv_2 \inv[2154]/_0_  (.A(\inv_in[2154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2155] ));
 sky130_fd_sc_hd__inv_2 \inv[2155]/_0_  (.A(\inv_in[2155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2156] ));
 sky130_fd_sc_hd__inv_2 \inv[2156]/_0_  (.A(\inv_in[2156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2157] ));
 sky130_fd_sc_hd__inv_2 \inv[2157]/_0_  (.A(\inv_in[2157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2158] ));
 sky130_fd_sc_hd__inv_2 \inv[2158]/_0_  (.A(\inv_in[2158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2159] ));
 sky130_fd_sc_hd__inv_2 \inv[2159]/_0_  (.A(\inv_in[2159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2160] ));
 sky130_fd_sc_hd__inv_2 \inv[215]/_0_  (.A(\inv_in[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[216] ));
 sky130_fd_sc_hd__inv_2 \inv[2160]/_0_  (.A(\inv_in[2160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2161] ));
 sky130_fd_sc_hd__inv_2 \inv[2161]/_0_  (.A(\inv_in[2161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2162] ));
 sky130_fd_sc_hd__inv_2 \inv[2162]/_0_  (.A(\inv_in[2162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2163] ));
 sky130_fd_sc_hd__inv_2 \inv[2163]/_0_  (.A(\inv_in[2163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2164] ));
 sky130_fd_sc_hd__inv_2 \inv[2164]/_0_  (.A(\inv_in[2164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2165] ));
 sky130_fd_sc_hd__inv_2 \inv[2165]/_0_  (.A(\inv_in[2165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2166] ));
 sky130_fd_sc_hd__inv_2 \inv[2166]/_0_  (.A(\inv_in[2166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2167] ));
 sky130_fd_sc_hd__inv_2 \inv[2167]/_0_  (.A(\inv_in[2167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2168] ));
 sky130_fd_sc_hd__inv_2 \inv[2168]/_0_  (.A(\inv_in[2168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2169] ));
 sky130_fd_sc_hd__inv_2 \inv[2169]/_0_  (.A(\inv_in[2169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2170] ));
 sky130_fd_sc_hd__inv_2 \inv[216]/_0_  (.A(\inv_in[216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[217] ));
 sky130_fd_sc_hd__inv_2 \inv[2170]/_0_  (.A(\inv_in[2170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2171] ));
 sky130_fd_sc_hd__inv_2 \inv[2171]/_0_  (.A(\inv_in[2171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2172] ));
 sky130_fd_sc_hd__inv_2 \inv[2172]/_0_  (.A(\inv_in[2172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2173] ));
 sky130_fd_sc_hd__inv_2 \inv[2173]/_0_  (.A(\inv_in[2173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2174] ));
 sky130_fd_sc_hd__inv_2 \inv[2174]/_0_  (.A(\inv_in[2174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2175] ));
 sky130_fd_sc_hd__inv_2 \inv[2175]/_0_  (.A(\inv_in[2175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2176] ));
 sky130_fd_sc_hd__inv_2 \inv[2176]/_0_  (.A(\inv_in[2176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2177] ));
 sky130_fd_sc_hd__inv_2 \inv[2177]/_0_  (.A(\inv_in[2177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2178] ));
 sky130_fd_sc_hd__inv_2 \inv[2178]/_0_  (.A(\inv_in[2178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2179] ));
 sky130_fd_sc_hd__inv_2 \inv[2179]/_0_  (.A(\inv_in[2179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2180] ));
 sky130_fd_sc_hd__inv_2 \inv[217]/_0_  (.A(\inv_in[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[218] ));
 sky130_fd_sc_hd__inv_2 \inv[2180]/_0_  (.A(\inv_in[2180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2181] ));
 sky130_fd_sc_hd__inv_2 \inv[2181]/_0_  (.A(\inv_in[2181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2182] ));
 sky130_fd_sc_hd__inv_2 \inv[2182]/_0_  (.A(\inv_in[2182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2183] ));
 sky130_fd_sc_hd__inv_2 \inv[2183]/_0_  (.A(\inv_in[2183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2184] ));
 sky130_fd_sc_hd__inv_2 \inv[2184]/_0_  (.A(\inv_in[2184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2185] ));
 sky130_fd_sc_hd__inv_2 \inv[2185]/_0_  (.A(\inv_in[2185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2186] ));
 sky130_fd_sc_hd__inv_2 \inv[2186]/_0_  (.A(\inv_in[2186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2187] ));
 sky130_fd_sc_hd__inv_2 \inv[2187]/_0_  (.A(\inv_in[2187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2188] ));
 sky130_fd_sc_hd__inv_2 \inv[2188]/_0_  (.A(\inv_in[2188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2189] ));
 sky130_fd_sc_hd__inv_2 \inv[2189]/_0_  (.A(\inv_in[2189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2190] ));
 sky130_fd_sc_hd__inv_2 \inv[218]/_0_  (.A(\inv_in[218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[219] ));
 sky130_fd_sc_hd__inv_2 \inv[2190]/_0_  (.A(\inv_in[2190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2191] ));
 sky130_fd_sc_hd__inv_2 \inv[2191]/_0_  (.A(\inv_in[2191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2192] ));
 sky130_fd_sc_hd__inv_2 \inv[2192]/_0_  (.A(\inv_in[2192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2193] ));
 sky130_fd_sc_hd__inv_2 \inv[2193]/_0_  (.A(\inv_in[2193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2194] ));
 sky130_fd_sc_hd__inv_2 \inv[2194]/_0_  (.A(\inv_in[2194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2195] ));
 sky130_fd_sc_hd__inv_2 \inv[2195]/_0_  (.A(\inv_in[2195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2196] ));
 sky130_fd_sc_hd__inv_2 \inv[2196]/_0_  (.A(\inv_in[2196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2197] ));
 sky130_fd_sc_hd__inv_2 \inv[2197]/_0_  (.A(\inv_in[2197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2198] ));
 sky130_fd_sc_hd__inv_2 \inv[2198]/_0_  (.A(\inv_in[2198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2199] ));
 sky130_fd_sc_hd__inv_2 \inv[2199]/_0_  (.A(\inv_in[2199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2200] ));
 sky130_fd_sc_hd__inv_2 \inv[219]/_0_  (.A(\inv_in[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[220] ));
 sky130_fd_sc_hd__inv_2 \inv[21]/_0_  (.A(\inv_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[22] ));
 sky130_fd_sc_hd__inv_2 \inv[2200]/_0_  (.A(\inv_in[2200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2201] ));
 sky130_fd_sc_hd__inv_2 \inv[2201]/_0_  (.A(\inv_in[2201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2202] ));
 sky130_fd_sc_hd__inv_2 \inv[2202]/_0_  (.A(\inv_in[2202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2203] ));
 sky130_fd_sc_hd__inv_2 \inv[2203]/_0_  (.A(\inv_in[2203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2204] ));
 sky130_fd_sc_hd__inv_2 \inv[2204]/_0_  (.A(\inv_in[2204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2205] ));
 sky130_fd_sc_hd__inv_2 \inv[2205]/_0_  (.A(\inv_in[2205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2206] ));
 sky130_fd_sc_hd__inv_2 \inv[2206]/_0_  (.A(\inv_in[2206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2207] ));
 sky130_fd_sc_hd__inv_2 \inv[2207]/_0_  (.A(\inv_in[2207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2208] ));
 sky130_fd_sc_hd__inv_2 \inv[2208]/_0_  (.A(\inv_in[2208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2209] ));
 sky130_fd_sc_hd__inv_2 \inv[2209]/_0_  (.A(\inv_in[2209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2210] ));
 sky130_fd_sc_hd__inv_2 \inv[220]/_0_  (.A(\inv_in[220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[221] ));
 sky130_fd_sc_hd__inv_2 \inv[2210]/_0_  (.A(\inv_in[2210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2211] ));
 sky130_fd_sc_hd__inv_2 \inv[2211]/_0_  (.A(\inv_in[2211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2212] ));
 sky130_fd_sc_hd__inv_2 \inv[2212]/_0_  (.A(\inv_in[2212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2213] ));
 sky130_fd_sc_hd__inv_2 \inv[2213]/_0_  (.A(\inv_in[2213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2214] ));
 sky130_fd_sc_hd__inv_2 \inv[2214]/_0_  (.A(\inv_in[2214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2215] ));
 sky130_fd_sc_hd__inv_2 \inv[2215]/_0_  (.A(\inv_in[2215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2216] ));
 sky130_fd_sc_hd__inv_2 \inv[2216]/_0_  (.A(\inv_in[2216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2217] ));
 sky130_fd_sc_hd__inv_2 \inv[2217]/_0_  (.A(\inv_in[2217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2218] ));
 sky130_fd_sc_hd__inv_2 \inv[2218]/_0_  (.A(\inv_in[2218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2219] ));
 sky130_fd_sc_hd__inv_2 \inv[2219]/_0_  (.A(\inv_in[2219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2220] ));
 sky130_fd_sc_hd__inv_2 \inv[221]/_0_  (.A(\inv_in[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[222] ));
 sky130_fd_sc_hd__inv_2 \inv[2220]/_0_  (.A(\inv_in[2220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2221] ));
 sky130_fd_sc_hd__inv_2 \inv[2221]/_0_  (.A(\inv_in[2221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2222] ));
 sky130_fd_sc_hd__inv_2 \inv[2222]/_0_  (.A(\inv_in[2222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2223] ));
 sky130_fd_sc_hd__inv_2 \inv[2223]/_0_  (.A(\inv_in[2223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2224] ));
 sky130_fd_sc_hd__inv_2 \inv[2224]/_0_  (.A(\inv_in[2224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2225] ));
 sky130_fd_sc_hd__inv_2 \inv[2225]/_0_  (.A(\inv_in[2225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2226] ));
 sky130_fd_sc_hd__inv_2 \inv[2226]/_0_  (.A(\inv_in[2226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2227] ));
 sky130_fd_sc_hd__inv_2 \inv[2227]/_0_  (.A(\inv_in[2227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2228] ));
 sky130_fd_sc_hd__inv_2 \inv[2228]/_0_  (.A(\inv_in[2228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2229] ));
 sky130_fd_sc_hd__inv_2 \inv[2229]/_0_  (.A(\inv_in[2229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2230] ));
 sky130_fd_sc_hd__inv_2 \inv[222]/_0_  (.A(\inv_in[222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[223] ));
 sky130_fd_sc_hd__inv_2 \inv[2230]/_0_  (.A(\inv_in[2230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2231] ));
 sky130_fd_sc_hd__inv_2 \inv[2231]/_0_  (.A(\inv_in[2231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2232] ));
 sky130_fd_sc_hd__inv_2 \inv[2232]/_0_  (.A(\inv_in[2232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2233] ));
 sky130_fd_sc_hd__inv_2 \inv[2233]/_0_  (.A(\inv_in[2233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2234] ));
 sky130_fd_sc_hd__inv_2 \inv[2234]/_0_  (.A(\inv_in[2234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2235] ));
 sky130_fd_sc_hd__inv_2 \inv[2235]/_0_  (.A(\inv_in[2235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2236] ));
 sky130_fd_sc_hd__inv_2 \inv[2236]/_0_  (.A(\inv_in[2236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2237] ));
 sky130_fd_sc_hd__inv_2 \inv[2237]/_0_  (.A(\inv_in[2237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2238] ));
 sky130_fd_sc_hd__inv_2 \inv[2238]/_0_  (.A(\inv_in[2238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2239] ));
 sky130_fd_sc_hd__inv_2 \inv[2239]/_0_  (.A(\inv_in[2239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2240] ));
 sky130_fd_sc_hd__inv_2 \inv[223]/_0_  (.A(\inv_in[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[224] ));
 sky130_fd_sc_hd__inv_2 \inv[2240]/_0_  (.A(\inv_in[2240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2241] ));
 sky130_fd_sc_hd__inv_2 \inv[2241]/_0_  (.A(\inv_in[2241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2242] ));
 sky130_fd_sc_hd__inv_2 \inv[2242]/_0_  (.A(\inv_in[2242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2243] ));
 sky130_fd_sc_hd__inv_2 \inv[2243]/_0_  (.A(\inv_in[2243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2244] ));
 sky130_fd_sc_hd__inv_2 \inv[2244]/_0_  (.A(\inv_in[2244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2245] ));
 sky130_fd_sc_hd__inv_2 \inv[2245]/_0_  (.A(\inv_in[2245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2246] ));
 sky130_fd_sc_hd__inv_2 \inv[2246]/_0_  (.A(\inv_in[2246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2247] ));
 sky130_fd_sc_hd__inv_2 \inv[2247]/_0_  (.A(\inv_in[2247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2248] ));
 sky130_fd_sc_hd__inv_2 \inv[2248]/_0_  (.A(\inv_in[2248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2249] ));
 sky130_fd_sc_hd__inv_2 \inv[2249]/_0_  (.A(\inv_in[2249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2250] ));
 sky130_fd_sc_hd__inv_2 \inv[224]/_0_  (.A(\inv_in[224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[225] ));
 sky130_fd_sc_hd__inv_2 \inv[2250]/_0_  (.A(\inv_in[2250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2251] ));
 sky130_fd_sc_hd__inv_2 \inv[2251]/_0_  (.A(\inv_in[2251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2252] ));
 sky130_fd_sc_hd__inv_2 \inv[2252]/_0_  (.A(\inv_in[2252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2253] ));
 sky130_fd_sc_hd__inv_2 \inv[2253]/_0_  (.A(\inv_in[2253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2254] ));
 sky130_fd_sc_hd__inv_2 \inv[2254]/_0_  (.A(\inv_in[2254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2255] ));
 sky130_fd_sc_hd__inv_2 \inv[2255]/_0_  (.A(\inv_in[2255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2256] ));
 sky130_fd_sc_hd__inv_2 \inv[2256]/_0_  (.A(\inv_in[2256] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2257] ));
 sky130_fd_sc_hd__inv_2 \inv[2257]/_0_  (.A(\inv_in[2257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2258] ));
 sky130_fd_sc_hd__inv_2 \inv[2258]/_0_  (.A(\inv_in[2258] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2259] ));
 sky130_fd_sc_hd__inv_2 \inv[2259]/_0_  (.A(\inv_in[2259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2260] ));
 sky130_fd_sc_hd__inv_2 \inv[225]/_0_  (.A(\inv_in[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[226] ));
 sky130_fd_sc_hd__inv_2 \inv[2260]/_0_  (.A(\inv_in[2260] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2261] ));
 sky130_fd_sc_hd__inv_2 \inv[2261]/_0_  (.A(\inv_in[2261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2262] ));
 sky130_fd_sc_hd__inv_2 \inv[2262]/_0_  (.A(\inv_in[2262] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2263] ));
 sky130_fd_sc_hd__inv_2 \inv[2263]/_0_  (.A(\inv_in[2263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2264] ));
 sky130_fd_sc_hd__inv_2 \inv[2264]/_0_  (.A(\inv_in[2264] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2265] ));
 sky130_fd_sc_hd__inv_2 \inv[2265]/_0_  (.A(\inv_in[2265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2266] ));
 sky130_fd_sc_hd__inv_2 \inv[2266]/_0_  (.A(\inv_in[2266] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2267] ));
 sky130_fd_sc_hd__inv_2 \inv[2267]/_0_  (.A(\inv_in[2267] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2268] ));
 sky130_fd_sc_hd__inv_2 \inv[2268]/_0_  (.A(\inv_in[2268] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2269] ));
 sky130_fd_sc_hd__inv_2 \inv[2269]/_0_  (.A(\inv_in[2269] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2270] ));
 sky130_fd_sc_hd__inv_2 \inv[226]/_0_  (.A(\inv_in[226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[227] ));
 sky130_fd_sc_hd__inv_2 \inv[2270]/_0_  (.A(\inv_in[2270] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2271] ));
 sky130_fd_sc_hd__inv_2 \inv[2271]/_0_  (.A(\inv_in[2271] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2272] ));
 sky130_fd_sc_hd__inv_2 \inv[2272]/_0_  (.A(\inv_in[2272] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2273] ));
 sky130_fd_sc_hd__inv_2 \inv[2273]/_0_  (.A(\inv_in[2273] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2274] ));
 sky130_fd_sc_hd__inv_2 \inv[2274]/_0_  (.A(\inv_in[2274] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2275] ));
 sky130_fd_sc_hd__inv_2 \inv[2275]/_0_  (.A(\inv_in[2275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2276] ));
 sky130_fd_sc_hd__inv_2 \inv[2276]/_0_  (.A(\inv_in[2276] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2277] ));
 sky130_fd_sc_hd__inv_2 \inv[2277]/_0_  (.A(\inv_in[2277] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2278] ));
 sky130_fd_sc_hd__inv_2 \inv[2278]/_0_  (.A(\inv_in[2278] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2279] ));
 sky130_fd_sc_hd__inv_2 \inv[2279]/_0_  (.A(\inv_in[2279] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2280] ));
 sky130_fd_sc_hd__inv_2 \inv[227]/_0_  (.A(\inv_in[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[228] ));
 sky130_fd_sc_hd__inv_2 \inv[2280]/_0_  (.A(\inv_in[2280] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2281] ));
 sky130_fd_sc_hd__inv_2 \inv[2281]/_0_  (.A(\inv_in[2281] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2282] ));
 sky130_fd_sc_hd__inv_2 \inv[2282]/_0_  (.A(\inv_in[2282] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2283] ));
 sky130_fd_sc_hd__inv_2 \inv[2283]/_0_  (.A(\inv_in[2283] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2284] ));
 sky130_fd_sc_hd__inv_2 \inv[2284]/_0_  (.A(\inv_in[2284] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2285] ));
 sky130_fd_sc_hd__inv_2 \inv[2285]/_0_  (.A(\inv_in[2285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2286] ));
 sky130_fd_sc_hd__inv_2 \inv[2286]/_0_  (.A(\inv_in[2286] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2287] ));
 sky130_fd_sc_hd__inv_2 \inv[2287]/_0_  (.A(\inv_in[2287] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2288] ));
 sky130_fd_sc_hd__inv_2 \inv[2288]/_0_  (.A(\inv_in[2288] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2289] ));
 sky130_fd_sc_hd__inv_2 \inv[2289]/_0_  (.A(\inv_in[2289] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2290] ));
 sky130_fd_sc_hd__inv_2 \inv[228]/_0_  (.A(\inv_in[228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[229] ));
 sky130_fd_sc_hd__inv_2 \inv[2290]/_0_  (.A(\inv_in[2290] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2291] ));
 sky130_fd_sc_hd__inv_2 \inv[2291]/_0_  (.A(\inv_in[2291] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2292] ));
 sky130_fd_sc_hd__inv_2 \inv[2292]/_0_  (.A(\inv_in[2292] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2293] ));
 sky130_fd_sc_hd__inv_2 \inv[2293]/_0_  (.A(\inv_in[2293] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2294] ));
 sky130_fd_sc_hd__inv_2 \inv[2294]/_0_  (.A(\inv_in[2294] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2295] ));
 sky130_fd_sc_hd__inv_2 \inv[2295]/_0_  (.A(\inv_in[2295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2296] ));
 sky130_fd_sc_hd__inv_2 \inv[2296]/_0_  (.A(\inv_in[2296] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2297] ));
 sky130_fd_sc_hd__inv_2 \inv[2297]/_0_  (.A(\inv_in[2297] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2298] ));
 sky130_fd_sc_hd__inv_2 \inv[2298]/_0_  (.A(\inv_in[2298] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2299] ));
 sky130_fd_sc_hd__inv_2 \inv[2299]/_0_  (.A(\inv_in[2299] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2300] ));
 sky130_fd_sc_hd__inv_2 \inv[229]/_0_  (.A(\inv_in[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[230] ));
 sky130_fd_sc_hd__inv_2 \inv[22]/_0_  (.A(\inv_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[23] ));
 sky130_fd_sc_hd__inv_2 \inv[2300]/_0_  (.A(\inv_in[2300] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2301] ));
 sky130_fd_sc_hd__inv_2 \inv[2301]/_0_  (.A(\inv_in[2301] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2302] ));
 sky130_fd_sc_hd__inv_2 \inv[2302]/_0_  (.A(\inv_in[2302] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2303] ));
 sky130_fd_sc_hd__inv_2 \inv[2303]/_0_  (.A(\inv_in[2303] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2304] ));
 sky130_fd_sc_hd__inv_2 \inv[2304]/_0_  (.A(\inv_in[2304] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2305] ));
 sky130_fd_sc_hd__inv_2 \inv[2305]/_0_  (.A(\inv_in[2305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2306] ));
 sky130_fd_sc_hd__inv_2 \inv[2306]/_0_  (.A(\inv_in[2306] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2307] ));
 sky130_fd_sc_hd__inv_2 \inv[2307]/_0_  (.A(\inv_in[2307] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2308] ));
 sky130_fd_sc_hd__inv_2 \inv[2308]/_0_  (.A(\inv_in[2308] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2309] ));
 sky130_fd_sc_hd__inv_2 \inv[2309]/_0_  (.A(\inv_in[2309] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2310] ));
 sky130_fd_sc_hd__inv_2 \inv[230]/_0_  (.A(\inv_in[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[231] ));
 sky130_fd_sc_hd__inv_2 \inv[2310]/_0_  (.A(\inv_in[2310] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2311] ));
 sky130_fd_sc_hd__inv_2 \inv[2311]/_0_  (.A(\inv_in[2311] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2312] ));
 sky130_fd_sc_hd__inv_2 \inv[2312]/_0_  (.A(\inv_in[2312] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2313] ));
 sky130_fd_sc_hd__inv_2 \inv[2313]/_0_  (.A(\inv_in[2313] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2314] ));
 sky130_fd_sc_hd__inv_2 \inv[2314]/_0_  (.A(\inv_in[2314] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2315] ));
 sky130_fd_sc_hd__inv_2 \inv[2315]/_0_  (.A(\inv_in[2315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2316] ));
 sky130_fd_sc_hd__inv_2 \inv[2316]/_0_  (.A(\inv_in[2316] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2317] ));
 sky130_fd_sc_hd__inv_2 \inv[2317]/_0_  (.A(\inv_in[2317] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2318] ));
 sky130_fd_sc_hd__inv_2 \inv[2318]/_0_  (.A(\inv_in[2318] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2319] ));
 sky130_fd_sc_hd__inv_2 \inv[2319]/_0_  (.A(\inv_in[2319] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2320] ));
 sky130_fd_sc_hd__inv_2 \inv[231]/_0_  (.A(\inv_in[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[232] ));
 sky130_fd_sc_hd__inv_2 \inv[2320]/_0_  (.A(\inv_in[2320] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2321] ));
 sky130_fd_sc_hd__inv_2 \inv[2321]/_0_  (.A(\inv_in[2321] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2322] ));
 sky130_fd_sc_hd__inv_2 \inv[2322]/_0_  (.A(\inv_in[2322] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2323] ));
 sky130_fd_sc_hd__inv_2 \inv[2323]/_0_  (.A(\inv_in[2323] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2324] ));
 sky130_fd_sc_hd__inv_2 \inv[2324]/_0_  (.A(\inv_in[2324] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2325] ));
 sky130_fd_sc_hd__inv_2 \inv[2325]/_0_  (.A(\inv_in[2325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2326] ));
 sky130_fd_sc_hd__inv_2 \inv[2326]/_0_  (.A(\inv_in[2326] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2327] ));
 sky130_fd_sc_hd__inv_2 \inv[2327]/_0_  (.A(\inv_in[2327] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2328] ));
 sky130_fd_sc_hd__inv_2 \inv[2328]/_0_  (.A(\inv_in[2328] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2329] ));
 sky130_fd_sc_hd__inv_2 \inv[2329]/_0_  (.A(\inv_in[2329] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2330] ));
 sky130_fd_sc_hd__inv_2 \inv[232]/_0_  (.A(\inv_in[232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[233] ));
 sky130_fd_sc_hd__inv_2 \inv[2330]/_0_  (.A(\inv_in[2330] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2331] ));
 sky130_fd_sc_hd__inv_2 \inv[2331]/_0_  (.A(\inv_in[2331] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2332] ));
 sky130_fd_sc_hd__inv_2 \inv[2332]/_0_  (.A(\inv_in[2332] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2333] ));
 sky130_fd_sc_hd__inv_2 \inv[2333]/_0_  (.A(\inv_in[2333] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2334] ));
 sky130_fd_sc_hd__inv_2 \inv[2334]/_0_  (.A(\inv_in[2334] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2335] ));
 sky130_fd_sc_hd__inv_2 \inv[2335]/_0_  (.A(\inv_in[2335] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2336] ));
 sky130_fd_sc_hd__inv_2 \inv[2336]/_0_  (.A(\inv_in[2336] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2337] ));
 sky130_fd_sc_hd__inv_2 \inv[2337]/_0_  (.A(\inv_in[2337] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2338] ));
 sky130_fd_sc_hd__inv_2 \inv[2338]/_0_  (.A(\inv_in[2338] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2339] ));
 sky130_fd_sc_hd__inv_2 \inv[2339]/_0_  (.A(\inv_in[2339] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2340] ));
 sky130_fd_sc_hd__inv_2 \inv[233]/_0_  (.A(\inv_in[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[234] ));
 sky130_fd_sc_hd__inv_2 \inv[2340]/_0_  (.A(\inv_in[2340] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2341] ));
 sky130_fd_sc_hd__inv_2 \inv[2341]/_0_  (.A(\inv_in[2341] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2342] ));
 sky130_fd_sc_hd__inv_2 \inv[2342]/_0_  (.A(\inv_in[2342] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2343] ));
 sky130_fd_sc_hd__inv_2 \inv[2343]/_0_  (.A(\inv_in[2343] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2344] ));
 sky130_fd_sc_hd__inv_2 \inv[2344]/_0_  (.A(\inv_in[2344] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2345] ));
 sky130_fd_sc_hd__inv_2 \inv[2345]/_0_  (.A(\inv_in[2345] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2346] ));
 sky130_fd_sc_hd__inv_2 \inv[2346]/_0_  (.A(\inv_in[2346] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2347] ));
 sky130_fd_sc_hd__inv_2 \inv[2347]/_0_  (.A(\inv_in[2347] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2348] ));
 sky130_fd_sc_hd__inv_2 \inv[2348]/_0_  (.A(\inv_in[2348] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2349] ));
 sky130_fd_sc_hd__inv_2 \inv[2349]/_0_  (.A(\inv_in[2349] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2350] ));
 sky130_fd_sc_hd__inv_2 \inv[234]/_0_  (.A(\inv_in[234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[235] ));
 sky130_fd_sc_hd__inv_2 \inv[2350]/_0_  (.A(\inv_in[2350] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2351] ));
 sky130_fd_sc_hd__inv_2 \inv[2351]/_0_  (.A(\inv_in[2351] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2352] ));
 sky130_fd_sc_hd__inv_2 \inv[2352]/_0_  (.A(\inv_in[2352] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2353] ));
 sky130_fd_sc_hd__inv_2 \inv[2353]/_0_  (.A(\inv_in[2353] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2354] ));
 sky130_fd_sc_hd__inv_2 \inv[2354]/_0_  (.A(\inv_in[2354] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2355] ));
 sky130_fd_sc_hd__inv_2 \inv[2355]/_0_  (.A(\inv_in[2355] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2356] ));
 sky130_fd_sc_hd__inv_2 \inv[2356]/_0_  (.A(\inv_in[2356] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2357] ));
 sky130_fd_sc_hd__inv_2 \inv[2357]/_0_  (.A(\inv_in[2357] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2358] ));
 sky130_fd_sc_hd__inv_2 \inv[2358]/_0_  (.A(\inv_in[2358] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2359] ));
 sky130_fd_sc_hd__inv_2 \inv[2359]/_0_  (.A(\inv_in[2359] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2360] ));
 sky130_fd_sc_hd__inv_2 \inv[235]/_0_  (.A(\inv_in[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[236] ));
 sky130_fd_sc_hd__inv_2 \inv[2360]/_0_  (.A(\inv_in[2360] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2361] ));
 sky130_fd_sc_hd__inv_2 \inv[2361]/_0_  (.A(\inv_in[2361] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2362] ));
 sky130_fd_sc_hd__inv_2 \inv[2362]/_0_  (.A(\inv_in[2362] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2363] ));
 sky130_fd_sc_hd__inv_2 \inv[2363]/_0_  (.A(\inv_in[2363] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2364] ));
 sky130_fd_sc_hd__inv_2 \inv[2364]/_0_  (.A(\inv_in[2364] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2365] ));
 sky130_fd_sc_hd__inv_2 \inv[2365]/_0_  (.A(\inv_in[2365] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2366] ));
 sky130_fd_sc_hd__inv_2 \inv[2366]/_0_  (.A(\inv_in[2366] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2367] ));
 sky130_fd_sc_hd__inv_2 \inv[2367]/_0_  (.A(\inv_in[2367] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2368] ));
 sky130_fd_sc_hd__inv_2 \inv[2368]/_0_  (.A(\inv_in[2368] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2369] ));
 sky130_fd_sc_hd__inv_2 \inv[2369]/_0_  (.A(\inv_in[2369] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2370] ));
 sky130_fd_sc_hd__inv_2 \inv[236]/_0_  (.A(\inv_in[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[237] ));
 sky130_fd_sc_hd__inv_2 \inv[2370]/_0_  (.A(\inv_in[2370] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2371] ));
 sky130_fd_sc_hd__inv_2 \inv[2371]/_0_  (.A(\inv_in[2371] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2372] ));
 sky130_fd_sc_hd__inv_2 \inv[2372]/_0_  (.A(\inv_in[2372] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2373] ));
 sky130_fd_sc_hd__inv_2 \inv[2373]/_0_  (.A(\inv_in[2373] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2374] ));
 sky130_fd_sc_hd__inv_2 \inv[2374]/_0_  (.A(\inv_in[2374] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2375] ));
 sky130_fd_sc_hd__inv_2 \inv[2375]/_0_  (.A(\inv_in[2375] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2376] ));
 sky130_fd_sc_hd__inv_2 \inv[2376]/_0_  (.A(\inv_in[2376] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2377] ));
 sky130_fd_sc_hd__inv_2 \inv[2377]/_0_  (.A(\inv_in[2377] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2378] ));
 sky130_fd_sc_hd__inv_2 \inv[2378]/_0_  (.A(\inv_in[2378] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2379] ));
 sky130_fd_sc_hd__inv_2 \inv[2379]/_0_  (.A(\inv_in[2379] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2380] ));
 sky130_fd_sc_hd__inv_2 \inv[237]/_0_  (.A(\inv_in[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[238] ));
 sky130_fd_sc_hd__inv_2 \inv[2380]/_0_  (.A(\inv_in[2380] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2381] ));
 sky130_fd_sc_hd__inv_2 \inv[2381]/_0_  (.A(\inv_in[2381] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2382] ));
 sky130_fd_sc_hd__inv_2 \inv[2382]/_0_  (.A(\inv_in[2382] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2383] ));
 sky130_fd_sc_hd__inv_2 \inv[2383]/_0_  (.A(\inv_in[2383] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2384] ));
 sky130_fd_sc_hd__inv_2 \inv[2384]/_0_  (.A(\inv_in[2384] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2385] ));
 sky130_fd_sc_hd__inv_2 \inv[2385]/_0_  (.A(\inv_in[2385] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2386] ));
 sky130_fd_sc_hd__inv_2 \inv[2386]/_0_  (.A(\inv_in[2386] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2387] ));
 sky130_fd_sc_hd__inv_2 \inv[2387]/_0_  (.A(\inv_in[2387] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2388] ));
 sky130_fd_sc_hd__inv_2 \inv[2388]/_0_  (.A(\inv_in[2388] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2389] ));
 sky130_fd_sc_hd__inv_2 \inv[2389]/_0_  (.A(\inv_in[2389] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2390] ));
 sky130_fd_sc_hd__inv_2 \inv[238]/_0_  (.A(\inv_in[238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[239] ));
 sky130_fd_sc_hd__inv_2 \inv[2390]/_0_  (.A(\inv_in[2390] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2391] ));
 sky130_fd_sc_hd__inv_2 \inv[2391]/_0_  (.A(\inv_in[2391] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2392] ));
 sky130_fd_sc_hd__inv_2 \inv[2392]/_0_  (.A(\inv_in[2392] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2393] ));
 sky130_fd_sc_hd__inv_2 \inv[2393]/_0_  (.A(\inv_in[2393] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2394] ));
 sky130_fd_sc_hd__inv_2 \inv[2394]/_0_  (.A(\inv_in[2394] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2395] ));
 sky130_fd_sc_hd__inv_2 \inv[2395]/_0_  (.A(\inv_in[2395] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2396] ));
 sky130_fd_sc_hd__inv_2 \inv[2396]/_0_  (.A(\inv_in[2396] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2397] ));
 sky130_fd_sc_hd__inv_2 \inv[2397]/_0_  (.A(\inv_in[2397] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2398] ));
 sky130_fd_sc_hd__inv_2 \inv[2398]/_0_  (.A(\inv_in[2398] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2399] ));
 sky130_fd_sc_hd__inv_2 \inv[2399]/_0_  (.A(\inv_in[2399] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2400] ));
 sky130_fd_sc_hd__inv_2 \inv[239]/_0_  (.A(\inv_in[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[240] ));
 sky130_fd_sc_hd__inv_2 \inv[23]/_0_  (.A(\inv_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[24] ));
 sky130_fd_sc_hd__inv_2 \inv[2400]/_0_  (.A(\inv_in[2400] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2401] ));
 sky130_fd_sc_hd__inv_2 \inv[2401]/_0_  (.A(\inv_in[2401] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2402] ));
 sky130_fd_sc_hd__inv_2 \inv[2402]/_0_  (.A(\inv_in[2402] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2403] ));
 sky130_fd_sc_hd__inv_2 \inv[2403]/_0_  (.A(\inv_in[2403] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2404] ));
 sky130_fd_sc_hd__inv_2 \inv[2404]/_0_  (.A(\inv_in[2404] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2405] ));
 sky130_fd_sc_hd__inv_2 \inv[2405]/_0_  (.A(\inv_in[2405] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2406] ));
 sky130_fd_sc_hd__inv_2 \inv[2406]/_0_  (.A(\inv_in[2406] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2407] ));
 sky130_fd_sc_hd__inv_2 \inv[2407]/_0_  (.A(\inv_in[2407] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2408] ));
 sky130_fd_sc_hd__inv_2 \inv[2408]/_0_  (.A(\inv_in[2408] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2409] ));
 sky130_fd_sc_hd__inv_2 \inv[2409]/_0_  (.A(\inv_in[2409] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2410] ));
 sky130_fd_sc_hd__inv_2 \inv[240]/_0_  (.A(\inv_in[240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[241] ));
 sky130_fd_sc_hd__inv_2 \inv[2410]/_0_  (.A(\inv_in[2410] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2411] ));
 sky130_fd_sc_hd__inv_2 \inv[2411]/_0_  (.A(\inv_in[2411] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2412] ));
 sky130_fd_sc_hd__inv_2 \inv[2412]/_0_  (.A(\inv_in[2412] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2413] ));
 sky130_fd_sc_hd__inv_2 \inv[2413]/_0_  (.A(\inv_in[2413] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2414] ));
 sky130_fd_sc_hd__inv_2 \inv[2414]/_0_  (.A(\inv_in[2414] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2415] ));
 sky130_fd_sc_hd__inv_2 \inv[2415]/_0_  (.A(\inv_in[2415] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2416] ));
 sky130_fd_sc_hd__inv_2 \inv[2416]/_0_  (.A(\inv_in[2416] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2417] ));
 sky130_fd_sc_hd__inv_2 \inv[2417]/_0_  (.A(\inv_in[2417] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2418] ));
 sky130_fd_sc_hd__inv_2 \inv[2418]/_0_  (.A(\inv_in[2418] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2419] ));
 sky130_fd_sc_hd__inv_2 \inv[2419]/_0_  (.A(\inv_in[2419] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2420] ));
 sky130_fd_sc_hd__inv_2 \inv[241]/_0_  (.A(\inv_in[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[242] ));
 sky130_fd_sc_hd__inv_2 \inv[2420]/_0_  (.A(\inv_in[2420] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2421] ));
 sky130_fd_sc_hd__inv_2 \inv[2421]/_0_  (.A(\inv_in[2421] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2422] ));
 sky130_fd_sc_hd__inv_2 \inv[2422]/_0_  (.A(\inv_in[2422] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2423] ));
 sky130_fd_sc_hd__inv_2 \inv[2423]/_0_  (.A(\inv_in[2423] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2424] ));
 sky130_fd_sc_hd__inv_2 \inv[2424]/_0_  (.A(\inv_in[2424] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2425] ));
 sky130_fd_sc_hd__inv_2 \inv[2425]/_0_  (.A(\inv_in[2425] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2426] ));
 sky130_fd_sc_hd__inv_2 \inv[2426]/_0_  (.A(\inv_in[2426] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2427] ));
 sky130_fd_sc_hd__inv_2 \inv[2427]/_0_  (.A(\inv_in[2427] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2428] ));
 sky130_fd_sc_hd__inv_2 \inv[2428]/_0_  (.A(\inv_in[2428] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2429] ));
 sky130_fd_sc_hd__inv_2 \inv[2429]/_0_  (.A(\inv_in[2429] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2430] ));
 sky130_fd_sc_hd__inv_2 \inv[242]/_0_  (.A(\inv_in[242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[243] ));
 sky130_fd_sc_hd__inv_2 \inv[2430]/_0_  (.A(\inv_in[2430] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2431] ));
 sky130_fd_sc_hd__inv_2 \inv[2431]/_0_  (.A(\inv_in[2431] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2432] ));
 sky130_fd_sc_hd__inv_2 \inv[2432]/_0_  (.A(\inv_in[2432] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2433] ));
 sky130_fd_sc_hd__inv_2 \inv[2433]/_0_  (.A(\inv_in[2433] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2434] ));
 sky130_fd_sc_hd__inv_2 \inv[2434]/_0_  (.A(\inv_in[2434] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2435] ));
 sky130_fd_sc_hd__inv_2 \inv[2435]/_0_  (.A(\inv_in[2435] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2436] ));
 sky130_fd_sc_hd__inv_2 \inv[2436]/_0_  (.A(\inv_in[2436] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2437] ));
 sky130_fd_sc_hd__inv_2 \inv[2437]/_0_  (.A(\inv_in[2437] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2438] ));
 sky130_fd_sc_hd__inv_2 \inv[2438]/_0_  (.A(\inv_in[2438] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2439] ));
 sky130_fd_sc_hd__inv_2 \inv[2439]/_0_  (.A(\inv_in[2439] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2440] ));
 sky130_fd_sc_hd__inv_2 \inv[243]/_0_  (.A(\inv_in[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[244] ));
 sky130_fd_sc_hd__inv_2 \inv[2440]/_0_  (.A(\inv_in[2440] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2441] ));
 sky130_fd_sc_hd__inv_2 \inv[2441]/_0_  (.A(\inv_in[2441] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2442] ));
 sky130_fd_sc_hd__inv_2 \inv[2442]/_0_  (.A(\inv_in[2442] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2443] ));
 sky130_fd_sc_hd__inv_2 \inv[2443]/_0_  (.A(\inv_in[2443] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2444] ));
 sky130_fd_sc_hd__inv_2 \inv[2444]/_0_  (.A(\inv_in[2444] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2445] ));
 sky130_fd_sc_hd__inv_2 \inv[2445]/_0_  (.A(\inv_in[2445] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2446] ));
 sky130_fd_sc_hd__inv_2 \inv[2446]/_0_  (.A(\inv_in[2446] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2447] ));
 sky130_fd_sc_hd__inv_2 \inv[2447]/_0_  (.A(\inv_in[2447] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2448] ));
 sky130_fd_sc_hd__inv_2 \inv[2448]/_0_  (.A(\inv_in[2448] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2449] ));
 sky130_fd_sc_hd__inv_2 \inv[2449]/_0_  (.A(\inv_in[2449] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2450] ));
 sky130_fd_sc_hd__inv_2 \inv[244]/_0_  (.A(\inv_in[244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[245] ));
 sky130_fd_sc_hd__inv_2 \inv[2450]/_0_  (.A(\inv_in[2450] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2451] ));
 sky130_fd_sc_hd__inv_2 \inv[2451]/_0_  (.A(\inv_in[2451] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2452] ));
 sky130_fd_sc_hd__inv_2 \inv[2452]/_0_  (.A(\inv_in[2452] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2453] ));
 sky130_fd_sc_hd__inv_2 \inv[2453]/_0_  (.A(\inv_in[2453] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2454] ));
 sky130_fd_sc_hd__inv_2 \inv[2454]/_0_  (.A(\inv_in[2454] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2455] ));
 sky130_fd_sc_hd__inv_2 \inv[2455]/_0_  (.A(\inv_in[2455] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2456] ));
 sky130_fd_sc_hd__inv_2 \inv[2456]/_0_  (.A(\inv_in[2456] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2457] ));
 sky130_fd_sc_hd__inv_2 \inv[2457]/_0_  (.A(\inv_in[2457] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2458] ));
 sky130_fd_sc_hd__inv_2 \inv[2458]/_0_  (.A(\inv_in[2458] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2459] ));
 sky130_fd_sc_hd__inv_2 \inv[2459]/_0_  (.A(\inv_in[2459] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2460] ));
 sky130_fd_sc_hd__inv_2 \inv[245]/_0_  (.A(\inv_in[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[246] ));
 sky130_fd_sc_hd__inv_2 \inv[2460]/_0_  (.A(\inv_in[2460] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2461] ));
 sky130_fd_sc_hd__inv_2 \inv[2461]/_0_  (.A(\inv_in[2461] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2462] ));
 sky130_fd_sc_hd__inv_2 \inv[2462]/_0_  (.A(\inv_in[2462] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2463] ));
 sky130_fd_sc_hd__inv_2 \inv[2463]/_0_  (.A(\inv_in[2463] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2464] ));
 sky130_fd_sc_hd__inv_2 \inv[2464]/_0_  (.A(\inv_in[2464] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2465] ));
 sky130_fd_sc_hd__inv_2 \inv[2465]/_0_  (.A(\inv_in[2465] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2466] ));
 sky130_fd_sc_hd__inv_2 \inv[2466]/_0_  (.A(\inv_in[2466] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2467] ));
 sky130_fd_sc_hd__inv_2 \inv[2467]/_0_  (.A(\inv_in[2467] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2468] ));
 sky130_fd_sc_hd__inv_2 \inv[2468]/_0_  (.A(\inv_in[2468] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2469] ));
 sky130_fd_sc_hd__inv_2 \inv[2469]/_0_  (.A(\inv_in[2469] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2470] ));
 sky130_fd_sc_hd__inv_2 \inv[246]/_0_  (.A(\inv_in[246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[247] ));
 sky130_fd_sc_hd__inv_2 \inv[2470]/_0_  (.A(\inv_in[2470] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2471] ));
 sky130_fd_sc_hd__inv_2 \inv[2471]/_0_  (.A(\inv_in[2471] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2472] ));
 sky130_fd_sc_hd__inv_2 \inv[2472]/_0_  (.A(\inv_in[2472] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2473] ));
 sky130_fd_sc_hd__inv_2 \inv[2473]/_0_  (.A(\inv_in[2473] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2474] ));
 sky130_fd_sc_hd__inv_2 \inv[2474]/_0_  (.A(\inv_in[2474] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2475] ));
 sky130_fd_sc_hd__inv_2 \inv[2475]/_0_  (.A(\inv_in[2475] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2476] ));
 sky130_fd_sc_hd__inv_2 \inv[2476]/_0_  (.A(\inv_in[2476] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2477] ));
 sky130_fd_sc_hd__inv_2 \inv[2477]/_0_  (.A(\inv_in[2477] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2478] ));
 sky130_fd_sc_hd__inv_2 \inv[2478]/_0_  (.A(\inv_in[2478] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2479] ));
 sky130_fd_sc_hd__inv_2 \inv[2479]/_0_  (.A(\inv_in[2479] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2480] ));
 sky130_fd_sc_hd__inv_2 \inv[247]/_0_  (.A(\inv_in[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[248] ));
 sky130_fd_sc_hd__inv_2 \inv[2480]/_0_  (.A(\inv_in[2480] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2481] ));
 sky130_fd_sc_hd__inv_2 \inv[2481]/_0_  (.A(\inv_in[2481] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2482] ));
 sky130_fd_sc_hd__inv_2 \inv[2482]/_0_  (.A(\inv_in[2482] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2483] ));
 sky130_fd_sc_hd__inv_2 \inv[2483]/_0_  (.A(\inv_in[2483] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2484] ));
 sky130_fd_sc_hd__inv_2 \inv[2484]/_0_  (.A(\inv_in[2484] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2485] ));
 sky130_fd_sc_hd__inv_2 \inv[2485]/_0_  (.A(\inv_in[2485] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2486] ));
 sky130_fd_sc_hd__inv_2 \inv[2486]/_0_  (.A(\inv_in[2486] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2487] ));
 sky130_fd_sc_hd__inv_2 \inv[2487]/_0_  (.A(\inv_in[2487] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2488] ));
 sky130_fd_sc_hd__inv_2 \inv[2488]/_0_  (.A(\inv_in[2488] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2489] ));
 sky130_fd_sc_hd__inv_2 \inv[2489]/_0_  (.A(\inv_in[2489] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2490] ));
 sky130_fd_sc_hd__inv_2 \inv[248]/_0_  (.A(\inv_in[248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[249] ));
 sky130_fd_sc_hd__inv_2 \inv[2490]/_0_  (.A(\inv_in[2490] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2491] ));
 sky130_fd_sc_hd__inv_2 \inv[2491]/_0_  (.A(\inv_in[2491] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2492] ));
 sky130_fd_sc_hd__inv_2 \inv[2492]/_0_  (.A(\inv_in[2492] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2493] ));
 sky130_fd_sc_hd__inv_2 \inv[2493]/_0_  (.A(\inv_in[2493] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2494] ));
 sky130_fd_sc_hd__inv_2 \inv[2494]/_0_  (.A(\inv_in[2494] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2495] ));
 sky130_fd_sc_hd__inv_2 \inv[2495]/_0_  (.A(\inv_in[2495] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2496] ));
 sky130_fd_sc_hd__inv_2 \inv[2496]/_0_  (.A(\inv_in[2496] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2497] ));
 sky130_fd_sc_hd__inv_2 \inv[2497]/_0_  (.A(\inv_in[2497] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2498] ));
 sky130_fd_sc_hd__inv_2 \inv[2498]/_0_  (.A(\inv_in[2498] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2499] ));
 sky130_fd_sc_hd__inv_2 \inv[2499]/_0_  (.A(\inv_in[2499] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2500] ));
 sky130_fd_sc_hd__inv_2 \inv[249]/_0_  (.A(\inv_in[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[250] ));
 sky130_fd_sc_hd__inv_2 \inv[24]/_0_  (.A(\inv_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[25] ));
 sky130_fd_sc_hd__inv_2 \inv[2500]/_0_  (.A(\inv_in[2500] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2501] ));
 sky130_fd_sc_hd__inv_2 \inv[2501]/_0_  (.A(\inv_in[2501] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2502] ));
 sky130_fd_sc_hd__inv_2 \inv[2502]/_0_  (.A(\inv_in[2502] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2503] ));
 sky130_fd_sc_hd__inv_2 \inv[2503]/_0_  (.A(\inv_in[2503] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2504] ));
 sky130_fd_sc_hd__inv_2 \inv[2504]/_0_  (.A(\inv_in[2504] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2505] ));
 sky130_fd_sc_hd__inv_2 \inv[2505]/_0_  (.A(\inv_in[2505] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2506] ));
 sky130_fd_sc_hd__inv_2 \inv[2506]/_0_  (.A(\inv_in[2506] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2507] ));
 sky130_fd_sc_hd__inv_2 \inv[2507]/_0_  (.A(\inv_in[2507] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2508] ));
 sky130_fd_sc_hd__inv_2 \inv[2508]/_0_  (.A(\inv_in[2508] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2509] ));
 sky130_fd_sc_hd__inv_2 \inv[2509]/_0_  (.A(\inv_in[2509] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2510] ));
 sky130_fd_sc_hd__inv_2 \inv[250]/_0_  (.A(\inv_in[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[251] ));
 sky130_fd_sc_hd__inv_2 \inv[2510]/_0_  (.A(\inv_in[2510] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2511] ));
 sky130_fd_sc_hd__inv_2 \inv[2511]/_0_  (.A(\inv_in[2511] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2512] ));
 sky130_fd_sc_hd__inv_2 \inv[2512]/_0_  (.A(\inv_in[2512] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2513] ));
 sky130_fd_sc_hd__inv_2 \inv[2513]/_0_  (.A(\inv_in[2513] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2514] ));
 sky130_fd_sc_hd__inv_2 \inv[2514]/_0_  (.A(\inv_in[2514] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2515] ));
 sky130_fd_sc_hd__inv_2 \inv[2515]/_0_  (.A(\inv_in[2515] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2516] ));
 sky130_fd_sc_hd__inv_2 \inv[2516]/_0_  (.A(\inv_in[2516] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2517] ));
 sky130_fd_sc_hd__inv_2 \inv[2517]/_0_  (.A(\inv_in[2517] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2518] ));
 sky130_fd_sc_hd__inv_2 \inv[2518]/_0_  (.A(\inv_in[2518] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2519] ));
 sky130_fd_sc_hd__inv_2 \inv[2519]/_0_  (.A(\inv_in[2519] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2520] ));
 sky130_fd_sc_hd__inv_2 \inv[251]/_0_  (.A(\inv_in[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[252] ));
 sky130_fd_sc_hd__inv_2 \inv[2520]/_0_  (.A(\inv_in[2520] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2521] ));
 sky130_fd_sc_hd__inv_2 \inv[2521]/_0_  (.A(\inv_in[2521] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2522] ));
 sky130_fd_sc_hd__inv_2 \inv[2522]/_0_  (.A(\inv_in[2522] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2523] ));
 sky130_fd_sc_hd__inv_2 \inv[2523]/_0_  (.A(\inv_in[2523] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2524] ));
 sky130_fd_sc_hd__inv_2 \inv[2524]/_0_  (.A(\inv_in[2524] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2525] ));
 sky130_fd_sc_hd__inv_2 \inv[2525]/_0_  (.A(\inv_in[2525] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2526] ));
 sky130_fd_sc_hd__inv_2 \inv[2526]/_0_  (.A(\inv_in[2526] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2527] ));
 sky130_fd_sc_hd__inv_2 \inv[2527]/_0_  (.A(\inv_in[2527] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2528] ));
 sky130_fd_sc_hd__inv_2 \inv[2528]/_0_  (.A(\inv_in[2528] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2529] ));
 sky130_fd_sc_hd__inv_2 \inv[2529]/_0_  (.A(\inv_in[2529] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2530] ));
 sky130_fd_sc_hd__inv_2 \inv[252]/_0_  (.A(\inv_in[252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[253] ));
 sky130_fd_sc_hd__inv_2 \inv[2530]/_0_  (.A(\inv_in[2530] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2531] ));
 sky130_fd_sc_hd__inv_2 \inv[2531]/_0_  (.A(\inv_in[2531] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2532] ));
 sky130_fd_sc_hd__inv_2 \inv[2532]/_0_  (.A(\inv_in[2532] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2533] ));
 sky130_fd_sc_hd__inv_2 \inv[2533]/_0_  (.A(\inv_in[2533] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2534] ));
 sky130_fd_sc_hd__inv_2 \inv[2534]/_0_  (.A(\inv_in[2534] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2535] ));
 sky130_fd_sc_hd__inv_2 \inv[2535]/_0_  (.A(\inv_in[2535] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2536] ));
 sky130_fd_sc_hd__inv_2 \inv[2536]/_0_  (.A(\inv_in[2536] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2537] ));
 sky130_fd_sc_hd__inv_2 \inv[2537]/_0_  (.A(\inv_in[2537] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2538] ));
 sky130_fd_sc_hd__inv_2 \inv[2538]/_0_  (.A(\inv_in[2538] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2539] ));
 sky130_fd_sc_hd__inv_2 \inv[2539]/_0_  (.A(\inv_in[2539] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2540] ));
 sky130_fd_sc_hd__inv_2 \inv[253]/_0_  (.A(\inv_in[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[254] ));
 sky130_fd_sc_hd__inv_2 \inv[2540]/_0_  (.A(\inv_in[2540] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2541] ));
 sky130_fd_sc_hd__inv_2 \inv[2541]/_0_  (.A(\inv_in[2541] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2542] ));
 sky130_fd_sc_hd__inv_2 \inv[2542]/_0_  (.A(\inv_in[2542] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2543] ));
 sky130_fd_sc_hd__inv_2 \inv[2543]/_0_  (.A(\inv_in[2543] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2544] ));
 sky130_fd_sc_hd__inv_2 \inv[2544]/_0_  (.A(\inv_in[2544] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2545] ));
 sky130_fd_sc_hd__inv_2 \inv[2545]/_0_  (.A(\inv_in[2545] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2546] ));
 sky130_fd_sc_hd__inv_2 \inv[2546]/_0_  (.A(\inv_in[2546] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2547] ));
 sky130_fd_sc_hd__inv_2 \inv[2547]/_0_  (.A(\inv_in[2547] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2548] ));
 sky130_fd_sc_hd__inv_2 \inv[2548]/_0_  (.A(\inv_in[2548] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2549] ));
 sky130_fd_sc_hd__inv_2 \inv[2549]/_0_  (.A(\inv_in[2549] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2550] ));
 sky130_fd_sc_hd__inv_2 \inv[254]/_0_  (.A(\inv_in[254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[255] ));
 sky130_fd_sc_hd__inv_2 \inv[2550]/_0_  (.A(\inv_in[2550] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2551] ));
 sky130_fd_sc_hd__inv_2 \inv[2551]/_0_  (.A(\inv_in[2551] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2552] ));
 sky130_fd_sc_hd__inv_2 \inv[2552]/_0_  (.A(\inv_in[2552] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2553] ));
 sky130_fd_sc_hd__inv_2 \inv[2553]/_0_  (.A(\inv_in[2553] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2554] ));
 sky130_fd_sc_hd__inv_2 \inv[2554]/_0_  (.A(\inv_in[2554] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2555] ));
 sky130_fd_sc_hd__inv_2 \inv[2555]/_0_  (.A(\inv_in[2555] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2556] ));
 sky130_fd_sc_hd__inv_2 \inv[2556]/_0_  (.A(\inv_in[2556] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2557] ));
 sky130_fd_sc_hd__inv_2 \inv[2557]/_0_  (.A(\inv_in[2557] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2558] ));
 sky130_fd_sc_hd__inv_2 \inv[2558]/_0_  (.A(\inv_in[2558] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2559] ));
 sky130_fd_sc_hd__inv_2 \inv[2559]/_0_  (.A(\inv_in[2559] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2560] ));
 sky130_fd_sc_hd__inv_2 \inv[255]/_0_  (.A(\inv_in[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[256] ));
 sky130_fd_sc_hd__inv_2 \inv[2560]/_0_  (.A(\inv_in[2560] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2561] ));
 sky130_fd_sc_hd__inv_2 \inv[2561]/_0_  (.A(\inv_in[2561] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2562] ));
 sky130_fd_sc_hd__inv_2 \inv[2562]/_0_  (.A(\inv_in[2562] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2563] ));
 sky130_fd_sc_hd__inv_2 \inv[2563]/_0_  (.A(\inv_in[2563] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2564] ));
 sky130_fd_sc_hd__inv_2 \inv[2564]/_0_  (.A(\inv_in[2564] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2565] ));
 sky130_fd_sc_hd__inv_2 \inv[2565]/_0_  (.A(\inv_in[2565] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2566] ));
 sky130_fd_sc_hd__inv_2 \inv[2566]/_0_  (.A(\inv_in[2566] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2567] ));
 sky130_fd_sc_hd__inv_2 \inv[2567]/_0_  (.A(\inv_in[2567] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2568] ));
 sky130_fd_sc_hd__inv_2 \inv[2568]/_0_  (.A(\inv_in[2568] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2569] ));
 sky130_fd_sc_hd__inv_2 \inv[2569]/_0_  (.A(\inv_in[2569] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2570] ));
 sky130_fd_sc_hd__inv_2 \inv[256]/_0_  (.A(\inv_in[256] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[257] ));
 sky130_fd_sc_hd__inv_2 \inv[2570]/_0_  (.A(\inv_in[2570] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2571] ));
 sky130_fd_sc_hd__inv_2 \inv[2571]/_0_  (.A(\inv_in[2571] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2572] ));
 sky130_fd_sc_hd__inv_2 \inv[2572]/_0_  (.A(\inv_in[2572] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2573] ));
 sky130_fd_sc_hd__inv_2 \inv[2573]/_0_  (.A(\inv_in[2573] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2574] ));
 sky130_fd_sc_hd__inv_2 \inv[2574]/_0_  (.A(\inv_in[2574] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2575] ));
 sky130_fd_sc_hd__inv_2 \inv[2575]/_0_  (.A(\inv_in[2575] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2576] ));
 sky130_fd_sc_hd__inv_2 \inv[2576]/_0_  (.A(\inv_in[2576] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2577] ));
 sky130_fd_sc_hd__inv_2 \inv[2577]/_0_  (.A(\inv_in[2577] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2578] ));
 sky130_fd_sc_hd__inv_2 \inv[2578]/_0_  (.A(\inv_in[2578] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2579] ));
 sky130_fd_sc_hd__inv_2 \inv[2579]/_0_  (.A(\inv_in[2579] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2580] ));
 sky130_fd_sc_hd__inv_2 \inv[257]/_0_  (.A(\inv_in[257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[258] ));
 sky130_fd_sc_hd__inv_2 \inv[2580]/_0_  (.A(\inv_in[2580] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2581] ));
 sky130_fd_sc_hd__inv_2 \inv[2581]/_0_  (.A(\inv_in[2581] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2582] ));
 sky130_fd_sc_hd__inv_2 \inv[2582]/_0_  (.A(\inv_in[2582] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2583] ));
 sky130_fd_sc_hd__inv_2 \inv[2583]/_0_  (.A(\inv_in[2583] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2584] ));
 sky130_fd_sc_hd__inv_2 \inv[2584]/_0_  (.A(\inv_in[2584] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2585] ));
 sky130_fd_sc_hd__inv_2 \inv[2585]/_0_  (.A(\inv_in[2585] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2586] ));
 sky130_fd_sc_hd__inv_2 \inv[2586]/_0_  (.A(\inv_in[2586] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2587] ));
 sky130_fd_sc_hd__inv_2 \inv[2587]/_0_  (.A(\inv_in[2587] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2588] ));
 sky130_fd_sc_hd__inv_2 \inv[2588]/_0_  (.A(\inv_in[2588] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2589] ));
 sky130_fd_sc_hd__inv_2 \inv[2589]/_0_  (.A(\inv_in[2589] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2590] ));
 sky130_fd_sc_hd__inv_2 \inv[258]/_0_  (.A(\inv_in[258] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[259] ));
 sky130_fd_sc_hd__inv_2 \inv[2590]/_0_  (.A(\inv_in[2590] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2591] ));
 sky130_fd_sc_hd__inv_2 \inv[2591]/_0_  (.A(\inv_in[2591] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2592] ));
 sky130_fd_sc_hd__inv_2 \inv[2592]/_0_  (.A(\inv_in[2592] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2593] ));
 sky130_fd_sc_hd__inv_2 \inv[2593]/_0_  (.A(\inv_in[2593] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2594] ));
 sky130_fd_sc_hd__inv_2 \inv[2594]/_0_  (.A(\inv_in[2594] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2595] ));
 sky130_fd_sc_hd__inv_2 \inv[2595]/_0_  (.A(\inv_in[2595] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2596] ));
 sky130_fd_sc_hd__inv_2 \inv[2596]/_0_  (.A(\inv_in[2596] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2597] ));
 sky130_fd_sc_hd__inv_2 \inv[2597]/_0_  (.A(\inv_in[2597] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2598] ));
 sky130_fd_sc_hd__inv_2 \inv[2598]/_0_  (.A(\inv_in[2598] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2599] ));
 sky130_fd_sc_hd__inv_2 \inv[2599]/_0_  (.A(\inv_in[2599] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2600] ));
 sky130_fd_sc_hd__inv_2 \inv[259]/_0_  (.A(\inv_in[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[260] ));
 sky130_fd_sc_hd__inv_2 \inv[25]/_0_  (.A(\inv_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[26] ));
 sky130_fd_sc_hd__inv_2 \inv[2600]/_0_  (.A(\inv_in[2600] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2601] ));
 sky130_fd_sc_hd__inv_2 \inv[2601]/_0_  (.A(\inv_in[2601] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2602] ));
 sky130_fd_sc_hd__inv_2 \inv[2602]/_0_  (.A(\inv_in[2602] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2603] ));
 sky130_fd_sc_hd__inv_2 \inv[2603]/_0_  (.A(\inv_in[2603] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2604] ));
 sky130_fd_sc_hd__inv_2 \inv[2604]/_0_  (.A(\inv_in[2604] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2605] ));
 sky130_fd_sc_hd__inv_2 \inv[2605]/_0_  (.A(\inv_in[2605] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2606] ));
 sky130_fd_sc_hd__inv_2 \inv[2606]/_0_  (.A(\inv_in[2606] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2607] ));
 sky130_fd_sc_hd__inv_2 \inv[2607]/_0_  (.A(\inv_in[2607] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2608] ));
 sky130_fd_sc_hd__inv_2 \inv[2608]/_0_  (.A(\inv_in[2608] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2609] ));
 sky130_fd_sc_hd__inv_2 \inv[2609]/_0_  (.A(\inv_in[2609] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2610] ));
 sky130_fd_sc_hd__inv_2 \inv[260]/_0_  (.A(\inv_in[260] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[261] ));
 sky130_fd_sc_hd__inv_2 \inv[2610]/_0_  (.A(\inv_in[2610] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2611] ));
 sky130_fd_sc_hd__inv_2 \inv[2611]/_0_  (.A(\inv_in[2611] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2612] ));
 sky130_fd_sc_hd__inv_2 \inv[2612]/_0_  (.A(\inv_in[2612] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2613] ));
 sky130_fd_sc_hd__inv_2 \inv[2613]/_0_  (.A(\inv_in[2613] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2614] ));
 sky130_fd_sc_hd__inv_2 \inv[2614]/_0_  (.A(\inv_in[2614] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2615] ));
 sky130_fd_sc_hd__inv_2 \inv[2615]/_0_  (.A(\inv_in[2615] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2616] ));
 sky130_fd_sc_hd__inv_2 \inv[2616]/_0_  (.A(\inv_in[2616] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2617] ));
 sky130_fd_sc_hd__inv_2 \inv[2617]/_0_  (.A(\inv_in[2617] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2618] ));
 sky130_fd_sc_hd__inv_2 \inv[2618]/_0_  (.A(\inv_in[2618] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2619] ));
 sky130_fd_sc_hd__inv_2 \inv[2619]/_0_  (.A(\inv_in[2619] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2620] ));
 sky130_fd_sc_hd__inv_2 \inv[261]/_0_  (.A(\inv_in[261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[262] ));
 sky130_fd_sc_hd__inv_2 \inv[2620]/_0_  (.A(\inv_in[2620] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2621] ));
 sky130_fd_sc_hd__inv_2 \inv[2621]/_0_  (.A(\inv_in[2621] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2622] ));
 sky130_fd_sc_hd__inv_2 \inv[2622]/_0_  (.A(\inv_in[2622] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2623] ));
 sky130_fd_sc_hd__inv_2 \inv[2623]/_0_  (.A(\inv_in[2623] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2624] ));
 sky130_fd_sc_hd__inv_2 \inv[2624]/_0_  (.A(\inv_in[2624] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2625] ));
 sky130_fd_sc_hd__inv_2 \inv[2625]/_0_  (.A(\inv_in[2625] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2626] ));
 sky130_fd_sc_hd__inv_2 \inv[2626]/_0_  (.A(\inv_in[2626] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2627] ));
 sky130_fd_sc_hd__inv_2 \inv[2627]/_0_  (.A(\inv_in[2627] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2628] ));
 sky130_fd_sc_hd__inv_2 \inv[2628]/_0_  (.A(\inv_in[2628] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2629] ));
 sky130_fd_sc_hd__inv_2 \inv[2629]/_0_  (.A(\inv_in[2629] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2630] ));
 sky130_fd_sc_hd__inv_2 \inv[262]/_0_  (.A(\inv_in[262] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[263] ));
 sky130_fd_sc_hd__inv_2 \inv[2630]/_0_  (.A(\inv_in[2630] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2631] ));
 sky130_fd_sc_hd__inv_2 \inv[2631]/_0_  (.A(\inv_in[2631] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2632] ));
 sky130_fd_sc_hd__inv_2 \inv[2632]/_0_  (.A(\inv_in[2632] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2633] ));
 sky130_fd_sc_hd__inv_2 \inv[2633]/_0_  (.A(\inv_in[2633] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2634] ));
 sky130_fd_sc_hd__inv_2 \inv[2634]/_0_  (.A(\inv_in[2634] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2635] ));
 sky130_fd_sc_hd__inv_2 \inv[2635]/_0_  (.A(\inv_in[2635] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2636] ));
 sky130_fd_sc_hd__inv_2 \inv[2636]/_0_  (.A(\inv_in[2636] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2637] ));
 sky130_fd_sc_hd__inv_2 \inv[2637]/_0_  (.A(\inv_in[2637] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2638] ));
 sky130_fd_sc_hd__inv_2 \inv[2638]/_0_  (.A(\inv_in[2638] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2639] ));
 sky130_fd_sc_hd__inv_2 \inv[2639]/_0_  (.A(\inv_in[2639] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2640] ));
 sky130_fd_sc_hd__inv_2 \inv[263]/_0_  (.A(\inv_in[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[264] ));
 sky130_fd_sc_hd__inv_2 \inv[2640]/_0_  (.A(\inv_in[2640] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2641] ));
 sky130_fd_sc_hd__inv_2 \inv[2641]/_0_  (.A(\inv_in[2641] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2642] ));
 sky130_fd_sc_hd__inv_2 \inv[2642]/_0_  (.A(\inv_in[2642] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2643] ));
 sky130_fd_sc_hd__inv_2 \inv[2643]/_0_  (.A(\inv_in[2643] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2644] ));
 sky130_fd_sc_hd__inv_2 \inv[2644]/_0_  (.A(\inv_in[2644] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2645] ));
 sky130_fd_sc_hd__inv_2 \inv[2645]/_0_  (.A(\inv_in[2645] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2646] ));
 sky130_fd_sc_hd__inv_2 \inv[2646]/_0_  (.A(\inv_in[2646] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2647] ));
 sky130_fd_sc_hd__inv_2 \inv[2647]/_0_  (.A(\inv_in[2647] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2648] ));
 sky130_fd_sc_hd__inv_2 \inv[2648]/_0_  (.A(\inv_in[2648] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2649] ));
 sky130_fd_sc_hd__inv_2 \inv[2649]/_0_  (.A(\inv_in[2649] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2650] ));
 sky130_fd_sc_hd__inv_2 \inv[264]/_0_  (.A(\inv_in[264] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[265] ));
 sky130_fd_sc_hd__inv_2 \inv[2650]/_0_  (.A(\inv_in[2650] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2651] ));
 sky130_fd_sc_hd__inv_2 \inv[2651]/_0_  (.A(\inv_in[2651] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2652] ));
 sky130_fd_sc_hd__inv_2 \inv[2652]/_0_  (.A(\inv_in[2652] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2653] ));
 sky130_fd_sc_hd__inv_2 \inv[2653]/_0_  (.A(\inv_in[2653] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2654] ));
 sky130_fd_sc_hd__inv_2 \inv[2654]/_0_  (.A(\inv_in[2654] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2655] ));
 sky130_fd_sc_hd__inv_2 \inv[2655]/_0_  (.A(\inv_in[2655] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2656] ));
 sky130_fd_sc_hd__inv_2 \inv[2656]/_0_  (.A(\inv_in[2656] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2657] ));
 sky130_fd_sc_hd__inv_2 \inv[2657]/_0_  (.A(\inv_in[2657] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2658] ));
 sky130_fd_sc_hd__inv_2 \inv[2658]/_0_  (.A(\inv_in[2658] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2659] ));
 sky130_fd_sc_hd__inv_2 \inv[2659]/_0_  (.A(\inv_in[2659] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2660] ));
 sky130_fd_sc_hd__inv_2 \inv[265]/_0_  (.A(\inv_in[265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[266] ));
 sky130_fd_sc_hd__inv_2 \inv[2660]/_0_  (.A(\inv_in[2660] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2661] ));
 sky130_fd_sc_hd__inv_2 \inv[2661]/_0_  (.A(\inv_in[2661] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2662] ));
 sky130_fd_sc_hd__inv_2 \inv[2662]/_0_  (.A(\inv_in[2662] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2663] ));
 sky130_fd_sc_hd__inv_2 \inv[2663]/_0_  (.A(\inv_in[2663] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2664] ));
 sky130_fd_sc_hd__inv_2 \inv[2664]/_0_  (.A(\inv_in[2664] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2665] ));
 sky130_fd_sc_hd__inv_2 \inv[2665]/_0_  (.A(\inv_in[2665] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2666] ));
 sky130_fd_sc_hd__inv_2 \inv[2666]/_0_  (.A(\inv_in[2666] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2667] ));
 sky130_fd_sc_hd__inv_2 \inv[2667]/_0_  (.A(\inv_in[2667] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2668] ));
 sky130_fd_sc_hd__inv_2 \inv[2668]/_0_  (.A(\inv_in[2668] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2669] ));
 sky130_fd_sc_hd__inv_2 \inv[2669]/_0_  (.A(\inv_in[2669] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2670] ));
 sky130_fd_sc_hd__inv_2 \inv[266]/_0_  (.A(\inv_in[266] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[267] ));
 sky130_fd_sc_hd__inv_2 \inv[2670]/_0_  (.A(\inv_in[2670] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2671] ));
 sky130_fd_sc_hd__inv_2 \inv[2671]/_0_  (.A(\inv_in[2671] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2672] ));
 sky130_fd_sc_hd__inv_2 \inv[2672]/_0_  (.A(\inv_in[2672] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2673] ));
 sky130_fd_sc_hd__inv_2 \inv[2673]/_0_  (.A(\inv_in[2673] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2674] ));
 sky130_fd_sc_hd__inv_2 \inv[2674]/_0_  (.A(\inv_in[2674] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2675] ));
 sky130_fd_sc_hd__inv_2 \inv[2675]/_0_  (.A(\inv_in[2675] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2676] ));
 sky130_fd_sc_hd__inv_2 \inv[2676]/_0_  (.A(\inv_in[2676] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2677] ));
 sky130_fd_sc_hd__inv_2 \inv[2677]/_0_  (.A(\inv_in[2677] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2678] ));
 sky130_fd_sc_hd__inv_2 \inv[2678]/_0_  (.A(\inv_in[2678] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2679] ));
 sky130_fd_sc_hd__inv_2 \inv[2679]/_0_  (.A(\inv_in[2679] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2680] ));
 sky130_fd_sc_hd__inv_2 \inv[267]/_0_  (.A(\inv_in[267] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[268] ));
 sky130_fd_sc_hd__inv_2 \inv[2680]/_0_  (.A(\inv_in[2680] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2681] ));
 sky130_fd_sc_hd__inv_2 \inv[2681]/_0_  (.A(\inv_in[2681] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2682] ));
 sky130_fd_sc_hd__inv_2 \inv[2682]/_0_  (.A(\inv_in[2682] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2683] ));
 sky130_fd_sc_hd__inv_2 \inv[2683]/_0_  (.A(\inv_in[2683] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2684] ));
 sky130_fd_sc_hd__inv_2 \inv[2684]/_0_  (.A(\inv_in[2684] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2685] ));
 sky130_fd_sc_hd__inv_2 \inv[2685]/_0_  (.A(\inv_in[2685] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2686] ));
 sky130_fd_sc_hd__inv_2 \inv[2686]/_0_  (.A(\inv_in[2686] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2687] ));
 sky130_fd_sc_hd__inv_2 \inv[2687]/_0_  (.A(\inv_in[2687] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2688] ));
 sky130_fd_sc_hd__inv_2 \inv[2688]/_0_  (.A(\inv_in[2688] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2689] ));
 sky130_fd_sc_hd__inv_2 \inv[2689]/_0_  (.A(\inv_in[2689] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2690] ));
 sky130_fd_sc_hd__inv_2 \inv[268]/_0_  (.A(\inv_in[268] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[269] ));
 sky130_fd_sc_hd__inv_2 \inv[2690]/_0_  (.A(\inv_in[2690] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2691] ));
 sky130_fd_sc_hd__inv_2 \inv[2691]/_0_  (.A(\inv_in[2691] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2692] ));
 sky130_fd_sc_hd__inv_2 \inv[2692]/_0_  (.A(\inv_in[2692] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2693] ));
 sky130_fd_sc_hd__inv_2 \inv[2693]/_0_  (.A(\inv_in[2693] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2694] ));
 sky130_fd_sc_hd__inv_2 \inv[2694]/_0_  (.A(\inv_in[2694] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2695] ));
 sky130_fd_sc_hd__inv_2 \inv[2695]/_0_  (.A(\inv_in[2695] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2696] ));
 sky130_fd_sc_hd__inv_2 \inv[2696]/_0_  (.A(\inv_in[2696] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2697] ));
 sky130_fd_sc_hd__inv_2 \inv[2697]/_0_  (.A(\inv_in[2697] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2698] ));
 sky130_fd_sc_hd__inv_2 \inv[2698]/_0_  (.A(\inv_in[2698] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2699] ));
 sky130_fd_sc_hd__inv_2 \inv[2699]/_0_  (.A(\inv_in[2699] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2700] ));
 sky130_fd_sc_hd__inv_2 \inv[269]/_0_  (.A(\inv_in[269] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[270] ));
 sky130_fd_sc_hd__inv_2 \inv[26]/_0_  (.A(\inv_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[27] ));
 sky130_fd_sc_hd__inv_2 \inv[2700]/_0_  (.A(\inv_in[2700] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2701] ));
 sky130_fd_sc_hd__inv_2 \inv[2701]/_0_  (.A(\inv_in[2701] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2702] ));
 sky130_fd_sc_hd__inv_2 \inv[2702]/_0_  (.A(\inv_in[2702] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2703] ));
 sky130_fd_sc_hd__inv_2 \inv[2703]/_0_  (.A(\inv_in[2703] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2704] ));
 sky130_fd_sc_hd__inv_2 \inv[2704]/_0_  (.A(\inv_in[2704] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2705] ));
 sky130_fd_sc_hd__inv_2 \inv[2705]/_0_  (.A(\inv_in[2705] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2706] ));
 sky130_fd_sc_hd__inv_2 \inv[2706]/_0_  (.A(\inv_in[2706] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2707] ));
 sky130_fd_sc_hd__inv_2 \inv[2707]/_0_  (.A(\inv_in[2707] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2708] ));
 sky130_fd_sc_hd__inv_2 \inv[2708]/_0_  (.A(\inv_in[2708] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2709] ));
 sky130_fd_sc_hd__inv_2 \inv[2709]/_0_  (.A(\inv_in[2709] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2710] ));
 sky130_fd_sc_hd__inv_2 \inv[270]/_0_  (.A(\inv_in[270] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[271] ));
 sky130_fd_sc_hd__inv_2 \inv[2710]/_0_  (.A(\inv_in[2710] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2711] ));
 sky130_fd_sc_hd__inv_2 \inv[2711]/_0_  (.A(\inv_in[2711] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2712] ));
 sky130_fd_sc_hd__inv_2 \inv[2712]/_0_  (.A(\inv_in[2712] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2713] ));
 sky130_fd_sc_hd__inv_2 \inv[2713]/_0_  (.A(\inv_in[2713] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2714] ));
 sky130_fd_sc_hd__inv_2 \inv[2714]/_0_  (.A(\inv_in[2714] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2715] ));
 sky130_fd_sc_hd__inv_2 \inv[2715]/_0_  (.A(\inv_in[2715] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2716] ));
 sky130_fd_sc_hd__inv_2 \inv[2716]/_0_  (.A(\inv_in[2716] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2717] ));
 sky130_fd_sc_hd__inv_2 \inv[2717]/_0_  (.A(\inv_in[2717] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2718] ));
 sky130_fd_sc_hd__inv_2 \inv[2718]/_0_  (.A(\inv_in[2718] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2719] ));
 sky130_fd_sc_hd__inv_2 \inv[2719]/_0_  (.A(\inv_in[2719] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2720] ));
 sky130_fd_sc_hd__inv_2 \inv[271]/_0_  (.A(\inv_in[271] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[272] ));
 sky130_fd_sc_hd__inv_2 \inv[2720]/_0_  (.A(\inv_in[2720] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2721] ));
 sky130_fd_sc_hd__inv_2 \inv[2721]/_0_  (.A(\inv_in[2721] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2722] ));
 sky130_fd_sc_hd__inv_2 \inv[2722]/_0_  (.A(\inv_in[2722] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2723] ));
 sky130_fd_sc_hd__inv_2 \inv[2723]/_0_  (.A(\inv_in[2723] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2724] ));
 sky130_fd_sc_hd__inv_2 \inv[2724]/_0_  (.A(\inv_in[2724] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2725] ));
 sky130_fd_sc_hd__inv_2 \inv[2725]/_0_  (.A(\inv_in[2725] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2726] ));
 sky130_fd_sc_hd__inv_2 \inv[2726]/_0_  (.A(\inv_in[2726] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2727] ));
 sky130_fd_sc_hd__inv_2 \inv[2727]/_0_  (.A(\inv_in[2727] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2728] ));
 sky130_fd_sc_hd__inv_2 \inv[2728]/_0_  (.A(\inv_in[2728] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2729] ));
 sky130_fd_sc_hd__inv_2 \inv[2729]/_0_  (.A(\inv_in[2729] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2730] ));
 sky130_fd_sc_hd__inv_2 \inv[272]/_0_  (.A(\inv_in[272] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[273] ));
 sky130_fd_sc_hd__inv_2 \inv[2730]/_0_  (.A(\inv_in[2730] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2731] ));
 sky130_fd_sc_hd__inv_2 \inv[2731]/_0_  (.A(\inv_in[2731] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2732] ));
 sky130_fd_sc_hd__inv_2 \inv[2732]/_0_  (.A(\inv_in[2732] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2733] ));
 sky130_fd_sc_hd__inv_2 \inv[2733]/_0_  (.A(\inv_in[2733] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2734] ));
 sky130_fd_sc_hd__inv_2 \inv[2734]/_0_  (.A(\inv_in[2734] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2735] ));
 sky130_fd_sc_hd__inv_2 \inv[2735]/_0_  (.A(\inv_in[2735] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2736] ));
 sky130_fd_sc_hd__inv_2 \inv[2736]/_0_  (.A(\inv_in[2736] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2737] ));
 sky130_fd_sc_hd__inv_2 \inv[2737]/_0_  (.A(\inv_in[2737] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2738] ));
 sky130_fd_sc_hd__inv_2 \inv[2738]/_0_  (.A(\inv_in[2738] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2739] ));
 sky130_fd_sc_hd__inv_2 \inv[2739]/_0_  (.A(\inv_in[2739] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2740] ));
 sky130_fd_sc_hd__inv_2 \inv[273]/_0_  (.A(\inv_in[273] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[274] ));
 sky130_fd_sc_hd__inv_2 \inv[2740]/_0_  (.A(\inv_in[2740] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2741] ));
 sky130_fd_sc_hd__inv_2 \inv[2741]/_0_  (.A(\inv_in[2741] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2742] ));
 sky130_fd_sc_hd__inv_2 \inv[2742]/_0_  (.A(\inv_in[2742] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2743] ));
 sky130_fd_sc_hd__inv_2 \inv[2743]/_0_  (.A(\inv_in[2743] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2744] ));
 sky130_fd_sc_hd__inv_2 \inv[2744]/_0_  (.A(\inv_in[2744] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2745] ));
 sky130_fd_sc_hd__inv_2 \inv[2745]/_0_  (.A(\inv_in[2745] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2746] ));
 sky130_fd_sc_hd__inv_2 \inv[2746]/_0_  (.A(\inv_in[2746] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2747] ));
 sky130_fd_sc_hd__inv_2 \inv[2747]/_0_  (.A(\inv_in[2747] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2748] ));
 sky130_fd_sc_hd__inv_2 \inv[2748]/_0_  (.A(\inv_in[2748] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2749] ));
 sky130_fd_sc_hd__inv_2 \inv[2749]/_0_  (.A(\inv_in[2749] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2750] ));
 sky130_fd_sc_hd__inv_2 \inv[274]/_0_  (.A(\inv_in[274] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[275] ));
 sky130_fd_sc_hd__inv_2 \inv[2750]/_0_  (.A(\inv_in[2750] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2751] ));
 sky130_fd_sc_hd__inv_2 \inv[2751]/_0_  (.A(\inv_in[2751] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2752] ));
 sky130_fd_sc_hd__inv_2 \inv[2752]/_0_  (.A(\inv_in[2752] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2753] ));
 sky130_fd_sc_hd__inv_2 \inv[2753]/_0_  (.A(\inv_in[2753] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2754] ));
 sky130_fd_sc_hd__inv_2 \inv[2754]/_0_  (.A(\inv_in[2754] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2755] ));
 sky130_fd_sc_hd__inv_2 \inv[2755]/_0_  (.A(\inv_in[2755] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2756] ));
 sky130_fd_sc_hd__inv_2 \inv[2756]/_0_  (.A(\inv_in[2756] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2757] ));
 sky130_fd_sc_hd__inv_2 \inv[2757]/_0_  (.A(\inv_in[2757] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2758] ));
 sky130_fd_sc_hd__inv_2 \inv[2758]/_0_  (.A(\inv_in[2758] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2759] ));
 sky130_fd_sc_hd__inv_2 \inv[2759]/_0_  (.A(\inv_in[2759] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2760] ));
 sky130_fd_sc_hd__inv_2 \inv[275]/_0_  (.A(\inv_in[275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[276] ));
 sky130_fd_sc_hd__inv_2 \inv[2760]/_0_  (.A(\inv_in[2760] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2761] ));
 sky130_fd_sc_hd__inv_2 \inv[2761]/_0_  (.A(\inv_in[2761] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2762] ));
 sky130_fd_sc_hd__inv_2 \inv[2762]/_0_  (.A(\inv_in[2762] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2763] ));
 sky130_fd_sc_hd__inv_2 \inv[2763]/_0_  (.A(\inv_in[2763] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2764] ));
 sky130_fd_sc_hd__inv_2 \inv[2764]/_0_  (.A(\inv_in[2764] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2765] ));
 sky130_fd_sc_hd__inv_2 \inv[2765]/_0_  (.A(\inv_in[2765] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2766] ));
 sky130_fd_sc_hd__inv_2 \inv[2766]/_0_  (.A(\inv_in[2766] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2767] ));
 sky130_fd_sc_hd__inv_2 \inv[2767]/_0_  (.A(\inv_in[2767] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2768] ));
 sky130_fd_sc_hd__inv_2 \inv[2768]/_0_  (.A(\inv_in[2768] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2769] ));
 sky130_fd_sc_hd__inv_2 \inv[2769]/_0_  (.A(\inv_in[2769] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2770] ));
 sky130_fd_sc_hd__inv_2 \inv[276]/_0_  (.A(\inv_in[276] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[277] ));
 sky130_fd_sc_hd__inv_2 \inv[2770]/_0_  (.A(\inv_in[2770] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2771] ));
 sky130_fd_sc_hd__inv_2 \inv[2771]/_0_  (.A(\inv_in[2771] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2772] ));
 sky130_fd_sc_hd__inv_2 \inv[2772]/_0_  (.A(\inv_in[2772] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2773] ));
 sky130_fd_sc_hd__inv_2 \inv[2773]/_0_  (.A(\inv_in[2773] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2774] ));
 sky130_fd_sc_hd__inv_2 \inv[2774]/_0_  (.A(\inv_in[2774] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2775] ));
 sky130_fd_sc_hd__inv_2 \inv[2775]/_0_  (.A(\inv_in[2775] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2776] ));
 sky130_fd_sc_hd__inv_2 \inv[2776]/_0_  (.A(\inv_in[2776] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2777] ));
 sky130_fd_sc_hd__inv_2 \inv[2777]/_0_  (.A(\inv_in[2777] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2778] ));
 sky130_fd_sc_hd__inv_2 \inv[2778]/_0_  (.A(\inv_in[2778] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2779] ));
 sky130_fd_sc_hd__inv_2 \inv[2779]/_0_  (.A(\inv_in[2779] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2780] ));
 sky130_fd_sc_hd__inv_2 \inv[277]/_0_  (.A(\inv_in[277] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[278] ));
 sky130_fd_sc_hd__inv_2 \inv[2780]/_0_  (.A(\inv_in[2780] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2781] ));
 sky130_fd_sc_hd__inv_2 \inv[2781]/_0_  (.A(\inv_in[2781] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2782] ));
 sky130_fd_sc_hd__inv_2 \inv[2782]/_0_  (.A(\inv_in[2782] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2783] ));
 sky130_fd_sc_hd__inv_2 \inv[2783]/_0_  (.A(\inv_in[2783] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2784] ));
 sky130_fd_sc_hd__inv_2 \inv[2784]/_0_  (.A(\inv_in[2784] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2785] ));
 sky130_fd_sc_hd__inv_2 \inv[2785]/_0_  (.A(\inv_in[2785] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2786] ));
 sky130_fd_sc_hd__inv_2 \inv[2786]/_0_  (.A(\inv_in[2786] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2787] ));
 sky130_fd_sc_hd__inv_2 \inv[2787]/_0_  (.A(\inv_in[2787] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2788] ));
 sky130_fd_sc_hd__inv_2 \inv[2788]/_0_  (.A(\inv_in[2788] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2789] ));
 sky130_fd_sc_hd__inv_2 \inv[2789]/_0_  (.A(\inv_in[2789] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2790] ));
 sky130_fd_sc_hd__inv_2 \inv[278]/_0_  (.A(\inv_in[278] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[279] ));
 sky130_fd_sc_hd__inv_2 \inv[2790]/_0_  (.A(\inv_in[2790] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2791] ));
 sky130_fd_sc_hd__inv_2 \inv[2791]/_0_  (.A(\inv_in[2791] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2792] ));
 sky130_fd_sc_hd__inv_2 \inv[2792]/_0_  (.A(\inv_in[2792] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2793] ));
 sky130_fd_sc_hd__inv_2 \inv[2793]/_0_  (.A(\inv_in[2793] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2794] ));
 sky130_fd_sc_hd__inv_2 \inv[2794]/_0_  (.A(\inv_in[2794] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2795] ));
 sky130_fd_sc_hd__inv_2 \inv[2795]/_0_  (.A(\inv_in[2795] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2796] ));
 sky130_fd_sc_hd__inv_2 \inv[2796]/_0_  (.A(\inv_in[2796] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2797] ));
 sky130_fd_sc_hd__inv_2 \inv[2797]/_0_  (.A(\inv_in[2797] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2798] ));
 sky130_fd_sc_hd__inv_2 \inv[2798]/_0_  (.A(\inv_in[2798] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2799] ));
 sky130_fd_sc_hd__inv_2 \inv[2799]/_0_  (.A(\inv_in[2799] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2800] ));
 sky130_fd_sc_hd__inv_2 \inv[279]/_0_  (.A(\inv_in[279] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[280] ));
 sky130_fd_sc_hd__inv_2 \inv[27]/_0_  (.A(\inv_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[28] ));
 sky130_fd_sc_hd__inv_2 \inv[2800]/_0_  (.A(\inv_in[2800] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2801] ));
 sky130_fd_sc_hd__inv_2 \inv[2801]/_0_  (.A(\inv_in[2801] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2802] ));
 sky130_fd_sc_hd__inv_2 \inv[2802]/_0_  (.A(\inv_in[2802] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2803] ));
 sky130_fd_sc_hd__inv_2 \inv[2803]/_0_  (.A(\inv_in[2803] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2804] ));
 sky130_fd_sc_hd__inv_2 \inv[2804]/_0_  (.A(\inv_in[2804] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2805] ));
 sky130_fd_sc_hd__inv_2 \inv[2805]/_0_  (.A(\inv_in[2805] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2806] ));
 sky130_fd_sc_hd__inv_2 \inv[2806]/_0_  (.A(\inv_in[2806] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2807] ));
 sky130_fd_sc_hd__inv_2 \inv[2807]/_0_  (.A(\inv_in[2807] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2808] ));
 sky130_fd_sc_hd__inv_2 \inv[2808]/_0_  (.A(\inv_in[2808] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2809] ));
 sky130_fd_sc_hd__inv_2 \inv[2809]/_0_  (.A(\inv_in[2809] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2810] ));
 sky130_fd_sc_hd__inv_2 \inv[280]/_0_  (.A(\inv_in[280] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[281] ));
 sky130_fd_sc_hd__inv_2 \inv[2810]/_0_  (.A(\inv_in[2810] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2811] ));
 sky130_fd_sc_hd__inv_2 \inv[2811]/_0_  (.A(\inv_in[2811] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2812] ));
 sky130_fd_sc_hd__inv_2 \inv[2812]/_0_  (.A(\inv_in[2812] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2813] ));
 sky130_fd_sc_hd__inv_2 \inv[2813]/_0_  (.A(\inv_in[2813] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2814] ));
 sky130_fd_sc_hd__inv_2 \inv[2814]/_0_  (.A(\inv_in[2814] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2815] ));
 sky130_fd_sc_hd__inv_2 \inv[2815]/_0_  (.A(\inv_in[2815] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2816] ));
 sky130_fd_sc_hd__inv_2 \inv[2816]/_0_  (.A(\inv_in[2816] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2817] ));
 sky130_fd_sc_hd__inv_2 \inv[2817]/_0_  (.A(\inv_in[2817] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2818] ));
 sky130_fd_sc_hd__inv_2 \inv[2818]/_0_  (.A(\inv_in[2818] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2819] ));
 sky130_fd_sc_hd__inv_2 \inv[2819]/_0_  (.A(\inv_in[2819] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2820] ));
 sky130_fd_sc_hd__inv_2 \inv[281]/_0_  (.A(\inv_in[281] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[282] ));
 sky130_fd_sc_hd__inv_2 \inv[2820]/_0_  (.A(\inv_in[2820] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2821] ));
 sky130_fd_sc_hd__inv_2 \inv[2821]/_0_  (.A(\inv_in[2821] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2822] ));
 sky130_fd_sc_hd__inv_2 \inv[2822]/_0_  (.A(\inv_in[2822] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2823] ));
 sky130_fd_sc_hd__inv_2 \inv[2823]/_0_  (.A(\inv_in[2823] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2824] ));
 sky130_fd_sc_hd__inv_2 \inv[2824]/_0_  (.A(\inv_in[2824] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2825] ));
 sky130_fd_sc_hd__inv_2 \inv[2825]/_0_  (.A(\inv_in[2825] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2826] ));
 sky130_fd_sc_hd__inv_2 \inv[2826]/_0_  (.A(\inv_in[2826] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2827] ));
 sky130_fd_sc_hd__inv_2 \inv[2827]/_0_  (.A(\inv_in[2827] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2828] ));
 sky130_fd_sc_hd__inv_2 \inv[2828]/_0_  (.A(\inv_in[2828] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2829] ));
 sky130_fd_sc_hd__inv_2 \inv[2829]/_0_  (.A(\inv_in[2829] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2830] ));
 sky130_fd_sc_hd__inv_2 \inv[282]/_0_  (.A(\inv_in[282] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[283] ));
 sky130_fd_sc_hd__inv_2 \inv[2830]/_0_  (.A(\inv_in[2830] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2831] ));
 sky130_fd_sc_hd__inv_2 \inv[2831]/_0_  (.A(\inv_in[2831] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2832] ));
 sky130_fd_sc_hd__inv_2 \inv[2832]/_0_  (.A(\inv_in[2832] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2833] ));
 sky130_fd_sc_hd__inv_2 \inv[2833]/_0_  (.A(\inv_in[2833] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2834] ));
 sky130_fd_sc_hd__inv_2 \inv[2834]/_0_  (.A(\inv_in[2834] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2835] ));
 sky130_fd_sc_hd__inv_2 \inv[2835]/_0_  (.A(\inv_in[2835] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2836] ));
 sky130_fd_sc_hd__inv_2 \inv[2836]/_0_  (.A(\inv_in[2836] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2837] ));
 sky130_fd_sc_hd__inv_2 \inv[2837]/_0_  (.A(\inv_in[2837] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2838] ));
 sky130_fd_sc_hd__inv_2 \inv[2838]/_0_  (.A(\inv_in[2838] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2839] ));
 sky130_fd_sc_hd__inv_2 \inv[2839]/_0_  (.A(\inv_in[2839] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2840] ));
 sky130_fd_sc_hd__inv_2 \inv[283]/_0_  (.A(\inv_in[283] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[284] ));
 sky130_fd_sc_hd__inv_2 \inv[2840]/_0_  (.A(\inv_in[2840] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2841] ));
 sky130_fd_sc_hd__inv_2 \inv[2841]/_0_  (.A(\inv_in[2841] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2842] ));
 sky130_fd_sc_hd__inv_2 \inv[2842]/_0_  (.A(\inv_in[2842] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2843] ));
 sky130_fd_sc_hd__inv_2 \inv[2843]/_0_  (.A(\inv_in[2843] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2844] ));
 sky130_fd_sc_hd__inv_2 \inv[2844]/_0_  (.A(\inv_in[2844] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2845] ));
 sky130_fd_sc_hd__inv_2 \inv[2845]/_0_  (.A(\inv_in[2845] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2846] ));
 sky130_fd_sc_hd__inv_2 \inv[2846]/_0_  (.A(\inv_in[2846] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2847] ));
 sky130_fd_sc_hd__inv_2 \inv[2847]/_0_  (.A(\inv_in[2847] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2848] ));
 sky130_fd_sc_hd__inv_2 \inv[2848]/_0_  (.A(\inv_in[2848] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2849] ));
 sky130_fd_sc_hd__inv_2 \inv[2849]/_0_  (.A(\inv_in[2849] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2850] ));
 sky130_fd_sc_hd__inv_2 \inv[284]/_0_  (.A(\inv_in[284] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[285] ));
 sky130_fd_sc_hd__inv_2 \inv[2850]/_0_  (.A(\inv_in[2850] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2851] ));
 sky130_fd_sc_hd__inv_2 \inv[2851]/_0_  (.A(\inv_in[2851] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2852] ));
 sky130_fd_sc_hd__inv_2 \inv[2852]/_0_  (.A(\inv_in[2852] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2853] ));
 sky130_fd_sc_hd__inv_2 \inv[2853]/_0_  (.A(\inv_in[2853] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2854] ));
 sky130_fd_sc_hd__inv_2 \inv[2854]/_0_  (.A(\inv_in[2854] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2855] ));
 sky130_fd_sc_hd__inv_2 \inv[2855]/_0_  (.A(\inv_in[2855] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2856] ));
 sky130_fd_sc_hd__inv_2 \inv[2856]/_0_  (.A(\inv_in[2856] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2857] ));
 sky130_fd_sc_hd__inv_2 \inv[2857]/_0_  (.A(\inv_in[2857] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2858] ));
 sky130_fd_sc_hd__inv_2 \inv[2858]/_0_  (.A(\inv_in[2858] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2859] ));
 sky130_fd_sc_hd__inv_2 \inv[2859]/_0_  (.A(\inv_in[2859] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2860] ));
 sky130_fd_sc_hd__inv_2 \inv[285]/_0_  (.A(\inv_in[285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[286] ));
 sky130_fd_sc_hd__inv_2 \inv[2860]/_0_  (.A(\inv_in[2860] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2861] ));
 sky130_fd_sc_hd__inv_2 \inv[2861]/_0_  (.A(\inv_in[2861] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2862] ));
 sky130_fd_sc_hd__inv_2 \inv[2862]/_0_  (.A(\inv_in[2862] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2863] ));
 sky130_fd_sc_hd__inv_2 \inv[2863]/_0_  (.A(\inv_in[2863] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2864] ));
 sky130_fd_sc_hd__inv_2 \inv[2864]/_0_  (.A(\inv_in[2864] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2865] ));
 sky130_fd_sc_hd__inv_2 \inv[2865]/_0_  (.A(\inv_in[2865] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2866] ));
 sky130_fd_sc_hd__inv_2 \inv[2866]/_0_  (.A(\inv_in[2866] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2867] ));
 sky130_fd_sc_hd__inv_2 \inv[2867]/_0_  (.A(\inv_in[2867] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2868] ));
 sky130_fd_sc_hd__inv_2 \inv[2868]/_0_  (.A(\inv_in[2868] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2869] ));
 sky130_fd_sc_hd__inv_2 \inv[2869]/_0_  (.A(\inv_in[2869] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2870] ));
 sky130_fd_sc_hd__inv_2 \inv[286]/_0_  (.A(\inv_in[286] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[287] ));
 sky130_fd_sc_hd__inv_2 \inv[2870]/_0_  (.A(\inv_in[2870] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2871] ));
 sky130_fd_sc_hd__inv_2 \inv[2871]/_0_  (.A(\inv_in[2871] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2872] ));
 sky130_fd_sc_hd__inv_2 \inv[2872]/_0_  (.A(\inv_in[2872] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2873] ));
 sky130_fd_sc_hd__inv_2 \inv[2873]/_0_  (.A(\inv_in[2873] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2874] ));
 sky130_fd_sc_hd__inv_2 \inv[2874]/_0_  (.A(\inv_in[2874] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2875] ));
 sky130_fd_sc_hd__inv_2 \inv[2875]/_0_  (.A(\inv_in[2875] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2876] ));
 sky130_fd_sc_hd__inv_2 \inv[2876]/_0_  (.A(\inv_in[2876] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2877] ));
 sky130_fd_sc_hd__inv_2 \inv[2877]/_0_  (.A(\inv_in[2877] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2878] ));
 sky130_fd_sc_hd__inv_2 \inv[2878]/_0_  (.A(\inv_in[2878] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2879] ));
 sky130_fd_sc_hd__inv_2 \inv[2879]/_0_  (.A(\inv_in[2879] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2880] ));
 sky130_fd_sc_hd__inv_2 \inv[287]/_0_  (.A(\inv_in[287] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[288] ));
 sky130_fd_sc_hd__inv_2 \inv[2880]/_0_  (.A(\inv_in[2880] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2881] ));
 sky130_fd_sc_hd__inv_2 \inv[2881]/_0_  (.A(\inv_in[2881] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2882] ));
 sky130_fd_sc_hd__inv_2 \inv[2882]/_0_  (.A(\inv_in[2882] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2883] ));
 sky130_fd_sc_hd__inv_2 \inv[2883]/_0_  (.A(\inv_in[2883] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2884] ));
 sky130_fd_sc_hd__inv_2 \inv[2884]/_0_  (.A(\inv_in[2884] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2885] ));
 sky130_fd_sc_hd__inv_2 \inv[2885]/_0_  (.A(\inv_in[2885] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2886] ));
 sky130_fd_sc_hd__inv_2 \inv[2886]/_0_  (.A(\inv_in[2886] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2887] ));
 sky130_fd_sc_hd__inv_2 \inv[2887]/_0_  (.A(\inv_in[2887] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2888] ));
 sky130_fd_sc_hd__inv_2 \inv[2888]/_0_  (.A(\inv_in[2888] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2889] ));
 sky130_fd_sc_hd__inv_2 \inv[2889]/_0_  (.A(\inv_in[2889] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2890] ));
 sky130_fd_sc_hd__inv_2 \inv[288]/_0_  (.A(\inv_in[288] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[289] ));
 sky130_fd_sc_hd__inv_2 \inv[2890]/_0_  (.A(\inv_in[2890] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2891] ));
 sky130_fd_sc_hd__inv_2 \inv[2891]/_0_  (.A(\inv_in[2891] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2892] ));
 sky130_fd_sc_hd__inv_2 \inv[2892]/_0_  (.A(\inv_in[2892] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2893] ));
 sky130_fd_sc_hd__inv_2 \inv[2893]/_0_  (.A(\inv_in[2893] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2894] ));
 sky130_fd_sc_hd__inv_2 \inv[2894]/_0_  (.A(\inv_in[2894] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2895] ));
 sky130_fd_sc_hd__inv_2 \inv[2895]/_0_  (.A(\inv_in[2895] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2896] ));
 sky130_fd_sc_hd__inv_2 \inv[2896]/_0_  (.A(\inv_in[2896] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2897] ));
 sky130_fd_sc_hd__inv_2 \inv[2897]/_0_  (.A(\inv_in[2897] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2898] ));
 sky130_fd_sc_hd__inv_2 \inv[2898]/_0_  (.A(\inv_in[2898] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2899] ));
 sky130_fd_sc_hd__inv_2 \inv[2899]/_0_  (.A(\inv_in[2899] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2900] ));
 sky130_fd_sc_hd__inv_2 \inv[289]/_0_  (.A(\inv_in[289] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[290] ));
 sky130_fd_sc_hd__inv_2 \inv[28]/_0_  (.A(\inv_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[29] ));
 sky130_fd_sc_hd__inv_2 \inv[2900]/_0_  (.A(\inv_in[2900] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2901] ));
 sky130_fd_sc_hd__inv_2 \inv[2901]/_0_  (.A(\inv_in[2901] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2902] ));
 sky130_fd_sc_hd__inv_2 \inv[2902]/_0_  (.A(\inv_in[2902] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2903] ));
 sky130_fd_sc_hd__inv_2 \inv[2903]/_0_  (.A(\inv_in[2903] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2904] ));
 sky130_fd_sc_hd__inv_2 \inv[2904]/_0_  (.A(\inv_in[2904] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2905] ));
 sky130_fd_sc_hd__inv_2 \inv[2905]/_0_  (.A(\inv_in[2905] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2906] ));
 sky130_fd_sc_hd__inv_2 \inv[2906]/_0_  (.A(\inv_in[2906] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2907] ));
 sky130_fd_sc_hd__inv_2 \inv[2907]/_0_  (.A(\inv_in[2907] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2908] ));
 sky130_fd_sc_hd__inv_2 \inv[2908]/_0_  (.A(\inv_in[2908] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2909] ));
 sky130_fd_sc_hd__inv_2 \inv[2909]/_0_  (.A(\inv_in[2909] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2910] ));
 sky130_fd_sc_hd__inv_2 \inv[290]/_0_  (.A(\inv_in[290] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[291] ));
 sky130_fd_sc_hd__inv_2 \inv[2910]/_0_  (.A(\inv_in[2910] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2911] ));
 sky130_fd_sc_hd__inv_2 \inv[2911]/_0_  (.A(\inv_in[2911] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2912] ));
 sky130_fd_sc_hd__inv_2 \inv[2912]/_0_  (.A(\inv_in[2912] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2913] ));
 sky130_fd_sc_hd__inv_2 \inv[2913]/_0_  (.A(\inv_in[2913] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2914] ));
 sky130_fd_sc_hd__inv_2 \inv[2914]/_0_  (.A(\inv_in[2914] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2915] ));
 sky130_fd_sc_hd__inv_2 \inv[2915]/_0_  (.A(\inv_in[2915] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2916] ));
 sky130_fd_sc_hd__inv_2 \inv[2916]/_0_  (.A(\inv_in[2916] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2917] ));
 sky130_fd_sc_hd__inv_2 \inv[2917]/_0_  (.A(\inv_in[2917] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2918] ));
 sky130_fd_sc_hd__inv_2 \inv[2918]/_0_  (.A(\inv_in[2918] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2919] ));
 sky130_fd_sc_hd__inv_2 \inv[2919]/_0_  (.A(\inv_in[2919] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2920] ));
 sky130_fd_sc_hd__inv_2 \inv[291]/_0_  (.A(\inv_in[291] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[292] ));
 sky130_fd_sc_hd__inv_2 \inv[2920]/_0_  (.A(\inv_in[2920] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2921] ));
 sky130_fd_sc_hd__inv_2 \inv[2921]/_0_  (.A(\inv_in[2921] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2922] ));
 sky130_fd_sc_hd__inv_2 \inv[2922]/_0_  (.A(\inv_in[2922] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2923] ));
 sky130_fd_sc_hd__inv_2 \inv[2923]/_0_  (.A(\inv_in[2923] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2924] ));
 sky130_fd_sc_hd__inv_2 \inv[2924]/_0_  (.A(\inv_in[2924] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2925] ));
 sky130_fd_sc_hd__inv_2 \inv[2925]/_0_  (.A(\inv_in[2925] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2926] ));
 sky130_fd_sc_hd__inv_2 \inv[2926]/_0_  (.A(\inv_in[2926] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2927] ));
 sky130_fd_sc_hd__inv_2 \inv[2927]/_0_  (.A(\inv_in[2927] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2928] ));
 sky130_fd_sc_hd__inv_2 \inv[2928]/_0_  (.A(\inv_in[2928] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2929] ));
 sky130_fd_sc_hd__inv_2 \inv[2929]/_0_  (.A(\inv_in[2929] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2930] ));
 sky130_fd_sc_hd__inv_2 \inv[292]/_0_  (.A(\inv_in[292] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[293] ));
 sky130_fd_sc_hd__inv_2 \inv[2930]/_0_  (.A(\inv_in[2930] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2931] ));
 sky130_fd_sc_hd__inv_2 \inv[2931]/_0_  (.A(\inv_in[2931] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2932] ));
 sky130_fd_sc_hd__inv_2 \inv[2932]/_0_  (.A(\inv_in[2932] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2933] ));
 sky130_fd_sc_hd__inv_2 \inv[2933]/_0_  (.A(\inv_in[2933] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2934] ));
 sky130_fd_sc_hd__inv_2 \inv[2934]/_0_  (.A(\inv_in[2934] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2935] ));
 sky130_fd_sc_hd__inv_2 \inv[2935]/_0_  (.A(\inv_in[2935] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2936] ));
 sky130_fd_sc_hd__inv_2 \inv[2936]/_0_  (.A(\inv_in[2936] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2937] ));
 sky130_fd_sc_hd__inv_2 \inv[2937]/_0_  (.A(\inv_in[2937] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2938] ));
 sky130_fd_sc_hd__inv_2 \inv[2938]/_0_  (.A(\inv_in[2938] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2939] ));
 sky130_fd_sc_hd__inv_2 \inv[2939]/_0_  (.A(\inv_in[2939] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2940] ));
 sky130_fd_sc_hd__inv_2 \inv[293]/_0_  (.A(\inv_in[293] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[294] ));
 sky130_fd_sc_hd__inv_2 \inv[2940]/_0_  (.A(\inv_in[2940] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2941] ));
 sky130_fd_sc_hd__inv_2 \inv[2941]/_0_  (.A(\inv_in[2941] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2942] ));
 sky130_fd_sc_hd__inv_2 \inv[2942]/_0_  (.A(\inv_in[2942] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2943] ));
 sky130_fd_sc_hd__inv_2 \inv[2943]/_0_  (.A(\inv_in[2943] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2944] ));
 sky130_fd_sc_hd__inv_2 \inv[2944]/_0_  (.A(\inv_in[2944] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2945] ));
 sky130_fd_sc_hd__inv_2 \inv[2945]/_0_  (.A(\inv_in[2945] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2946] ));
 sky130_fd_sc_hd__inv_2 \inv[2946]/_0_  (.A(\inv_in[2946] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2947] ));
 sky130_fd_sc_hd__inv_2 \inv[2947]/_0_  (.A(\inv_in[2947] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2948] ));
 sky130_fd_sc_hd__inv_2 \inv[2948]/_0_  (.A(\inv_in[2948] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2949] ));
 sky130_fd_sc_hd__inv_2 \inv[2949]/_0_  (.A(\inv_in[2949] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2950] ));
 sky130_fd_sc_hd__inv_2 \inv[294]/_0_  (.A(\inv_in[294] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[295] ));
 sky130_fd_sc_hd__inv_2 \inv[2950]/_0_  (.A(\inv_in[2950] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2951] ));
 sky130_fd_sc_hd__inv_2 \inv[2951]/_0_  (.A(\inv_in[2951] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2952] ));
 sky130_fd_sc_hd__inv_2 \inv[2952]/_0_  (.A(\inv_in[2952] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2953] ));
 sky130_fd_sc_hd__inv_2 \inv[2953]/_0_  (.A(\inv_in[2953] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2954] ));
 sky130_fd_sc_hd__inv_2 \inv[2954]/_0_  (.A(\inv_in[2954] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2955] ));
 sky130_fd_sc_hd__inv_2 \inv[2955]/_0_  (.A(\inv_in[2955] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2956] ));
 sky130_fd_sc_hd__inv_2 \inv[2956]/_0_  (.A(\inv_in[2956] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2957] ));
 sky130_fd_sc_hd__inv_2 \inv[2957]/_0_  (.A(\inv_in[2957] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2958] ));
 sky130_fd_sc_hd__inv_2 \inv[2958]/_0_  (.A(\inv_in[2958] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2959] ));
 sky130_fd_sc_hd__inv_2 \inv[2959]/_0_  (.A(\inv_in[2959] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2960] ));
 sky130_fd_sc_hd__inv_2 \inv[295]/_0_  (.A(\inv_in[295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[296] ));
 sky130_fd_sc_hd__inv_2 \inv[2960]/_0_  (.A(\inv_in[2960] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2961] ));
 sky130_fd_sc_hd__inv_2 \inv[2961]/_0_  (.A(\inv_in[2961] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2962] ));
 sky130_fd_sc_hd__inv_2 \inv[2962]/_0_  (.A(\inv_in[2962] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2963] ));
 sky130_fd_sc_hd__inv_2 \inv[2963]/_0_  (.A(\inv_in[2963] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2964] ));
 sky130_fd_sc_hd__inv_2 \inv[2964]/_0_  (.A(\inv_in[2964] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2965] ));
 sky130_fd_sc_hd__inv_2 \inv[2965]/_0_  (.A(\inv_in[2965] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2966] ));
 sky130_fd_sc_hd__inv_2 \inv[2966]/_0_  (.A(\inv_in[2966] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2967] ));
 sky130_fd_sc_hd__inv_2 \inv[2967]/_0_  (.A(\inv_in[2967] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2968] ));
 sky130_fd_sc_hd__inv_2 \inv[2968]/_0_  (.A(\inv_in[2968] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2969] ));
 sky130_fd_sc_hd__inv_2 \inv[2969]/_0_  (.A(\inv_in[2969] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2970] ));
 sky130_fd_sc_hd__inv_2 \inv[296]/_0_  (.A(\inv_in[296] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[297] ));
 sky130_fd_sc_hd__inv_2 \inv[2970]/_0_  (.A(\inv_in[2970] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2971] ));
 sky130_fd_sc_hd__inv_2 \inv[2971]/_0_  (.A(\inv_in[2971] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2972] ));
 sky130_fd_sc_hd__inv_2 \inv[2972]/_0_  (.A(\inv_in[2972] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2973] ));
 sky130_fd_sc_hd__inv_2 \inv[2973]/_0_  (.A(\inv_in[2973] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2974] ));
 sky130_fd_sc_hd__inv_2 \inv[2974]/_0_  (.A(\inv_in[2974] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2975] ));
 sky130_fd_sc_hd__inv_2 \inv[2975]/_0_  (.A(\inv_in[2975] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2976] ));
 sky130_fd_sc_hd__inv_2 \inv[2976]/_0_  (.A(\inv_in[2976] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2977] ));
 sky130_fd_sc_hd__inv_2 \inv[2977]/_0_  (.A(\inv_in[2977] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2978] ));
 sky130_fd_sc_hd__inv_2 \inv[2978]/_0_  (.A(\inv_in[2978] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2979] ));
 sky130_fd_sc_hd__inv_2 \inv[2979]/_0_  (.A(\inv_in[2979] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2980] ));
 sky130_fd_sc_hd__inv_2 \inv[297]/_0_  (.A(\inv_in[297] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[298] ));
 sky130_fd_sc_hd__inv_2 \inv[2980]/_0_  (.A(\inv_in[2980] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2981] ));
 sky130_fd_sc_hd__inv_2 \inv[2981]/_0_  (.A(\inv_in[2981] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2982] ));
 sky130_fd_sc_hd__inv_2 \inv[2982]/_0_  (.A(\inv_in[2982] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2983] ));
 sky130_fd_sc_hd__inv_2 \inv[2983]/_0_  (.A(\inv_in[2983] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2984] ));
 sky130_fd_sc_hd__inv_2 \inv[2984]/_0_  (.A(\inv_in[2984] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2985] ));
 sky130_fd_sc_hd__inv_2 \inv[2985]/_0_  (.A(\inv_in[2985] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2986] ));
 sky130_fd_sc_hd__inv_2 \inv[2986]/_0_  (.A(\inv_in[2986] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2987] ));
 sky130_fd_sc_hd__inv_2 \inv[2987]/_0_  (.A(\inv_in[2987] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2988] ));
 sky130_fd_sc_hd__inv_2 \inv[2988]/_0_  (.A(\inv_in[2988] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2989] ));
 sky130_fd_sc_hd__inv_2 \inv[2989]/_0_  (.A(\inv_in[2989] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2990] ));
 sky130_fd_sc_hd__inv_2 \inv[298]/_0_  (.A(\inv_in[298] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[299] ));
 sky130_fd_sc_hd__inv_2 \inv[2990]/_0_  (.A(\inv_in[2990] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2991] ));
 sky130_fd_sc_hd__inv_2 \inv[2991]/_0_  (.A(\inv_in[2991] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2992] ));
 sky130_fd_sc_hd__inv_2 \inv[2992]/_0_  (.A(\inv_in[2992] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2993] ));
 sky130_fd_sc_hd__inv_2 \inv[2993]/_0_  (.A(\inv_in[2993] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2994] ));
 sky130_fd_sc_hd__inv_2 \inv[2994]/_0_  (.A(\inv_in[2994] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2995] ));
 sky130_fd_sc_hd__inv_2 \inv[2995]/_0_  (.A(\inv_in[2995] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2996] ));
 sky130_fd_sc_hd__inv_2 \inv[2996]/_0_  (.A(\inv_in[2996] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2997] ));
 sky130_fd_sc_hd__inv_2 \inv[2997]/_0_  (.A(\inv_in[2997] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2998] ));
 sky130_fd_sc_hd__inv_2 \inv[2998]/_0_  (.A(\inv_in[2998] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[2999] ));
 sky130_fd_sc_hd__inv_2 \inv[2999]/_0_  (.A(\inv_in[2999] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3000] ));
 sky130_fd_sc_hd__inv_2 \inv[299]/_0_  (.A(\inv_in[299] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[300] ));
 sky130_fd_sc_hd__inv_2 \inv[29]/_0_  (.A(\inv_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[30] ));
 sky130_fd_sc_hd__inv_2 \inv[2]/_0_  (.A(\inv_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3] ));
 sky130_fd_sc_hd__inv_2 \inv[3000]/_0_  (.A(\inv_in[3000] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3001] ));
 sky130_fd_sc_hd__inv_2 \inv[3001]/_0_  (.A(\inv_in[3001] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3002] ));
 sky130_fd_sc_hd__inv_2 \inv[3002]/_0_  (.A(\inv_in[3002] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3003] ));
 sky130_fd_sc_hd__inv_2 \inv[3003]/_0_  (.A(\inv_in[3003] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3004] ));
 sky130_fd_sc_hd__inv_2 \inv[3004]/_0_  (.A(\inv_in[3004] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3005] ));
 sky130_fd_sc_hd__inv_2 \inv[3005]/_0_  (.A(\inv_in[3005] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3006] ));
 sky130_fd_sc_hd__inv_2 \inv[3006]/_0_  (.A(\inv_in[3006] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3007] ));
 sky130_fd_sc_hd__inv_2 \inv[3007]/_0_  (.A(\inv_in[3007] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3008] ));
 sky130_fd_sc_hd__inv_2 \inv[3008]/_0_  (.A(\inv_in[3008] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3009] ));
 sky130_fd_sc_hd__inv_2 \inv[3009]/_0_  (.A(\inv_in[3009] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3010] ));
 sky130_fd_sc_hd__inv_2 \inv[300]/_0_  (.A(\inv_in[300] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[301] ));
 sky130_fd_sc_hd__inv_2 \inv[3010]/_0_  (.A(\inv_in[3010] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3011] ));
 sky130_fd_sc_hd__inv_2 \inv[3011]/_0_  (.A(\inv_in[3011] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3012] ));
 sky130_fd_sc_hd__inv_2 \inv[3012]/_0_  (.A(\inv_in[3012] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3013] ));
 sky130_fd_sc_hd__inv_2 \inv[3013]/_0_  (.A(\inv_in[3013] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3014] ));
 sky130_fd_sc_hd__inv_2 \inv[3014]/_0_  (.A(\inv_in[3014] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3015] ));
 sky130_fd_sc_hd__inv_2 \inv[3015]/_0_  (.A(\inv_in[3015] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3016] ));
 sky130_fd_sc_hd__inv_2 \inv[3016]/_0_  (.A(\inv_in[3016] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3017] ));
 sky130_fd_sc_hd__inv_2 \inv[3017]/_0_  (.A(\inv_in[3017] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3018] ));
 sky130_fd_sc_hd__inv_2 \inv[3018]/_0_  (.A(\inv_in[3018] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3019] ));
 sky130_fd_sc_hd__inv_2 \inv[3019]/_0_  (.A(\inv_in[3019] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3020] ));
 sky130_fd_sc_hd__inv_2 \inv[301]/_0_  (.A(\inv_in[301] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[302] ));
 sky130_fd_sc_hd__inv_2 \inv[3020]/_0_  (.A(\inv_in[3020] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3021] ));
 sky130_fd_sc_hd__inv_2 \inv[3021]/_0_  (.A(\inv_in[3021] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3022] ));
 sky130_fd_sc_hd__inv_2 \inv[3022]/_0_  (.A(\inv_in[3022] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3023] ));
 sky130_fd_sc_hd__inv_2 \inv[3023]/_0_  (.A(\inv_in[3023] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3024] ));
 sky130_fd_sc_hd__inv_2 \inv[3024]/_0_  (.A(\inv_in[3024] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3025] ));
 sky130_fd_sc_hd__inv_2 \inv[3025]/_0_  (.A(\inv_in[3025] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3026] ));
 sky130_fd_sc_hd__inv_2 \inv[3026]/_0_  (.A(\inv_in[3026] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3027] ));
 sky130_fd_sc_hd__inv_2 \inv[3027]/_0_  (.A(\inv_in[3027] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3028] ));
 sky130_fd_sc_hd__inv_2 \inv[3028]/_0_  (.A(\inv_in[3028] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3029] ));
 sky130_fd_sc_hd__inv_2 \inv[3029]/_0_  (.A(\inv_in[3029] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3030] ));
 sky130_fd_sc_hd__inv_2 \inv[302]/_0_  (.A(\inv_in[302] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[303] ));
 sky130_fd_sc_hd__inv_2 \inv[3030]/_0_  (.A(\inv_in[3030] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3031] ));
 sky130_fd_sc_hd__inv_2 \inv[3031]/_0_  (.A(\inv_in[3031] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3032] ));
 sky130_fd_sc_hd__inv_2 \inv[3032]/_0_  (.A(\inv_in[3032] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3033] ));
 sky130_fd_sc_hd__inv_2 \inv[3033]/_0_  (.A(\inv_in[3033] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3034] ));
 sky130_fd_sc_hd__inv_2 \inv[3034]/_0_  (.A(\inv_in[3034] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3035] ));
 sky130_fd_sc_hd__inv_2 \inv[3035]/_0_  (.A(\inv_in[3035] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3036] ));
 sky130_fd_sc_hd__inv_2 \inv[3036]/_0_  (.A(\inv_in[3036] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3037] ));
 sky130_fd_sc_hd__inv_2 \inv[3037]/_0_  (.A(\inv_in[3037] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3038] ));
 sky130_fd_sc_hd__inv_2 \inv[3038]/_0_  (.A(\inv_in[3038] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3039] ));
 sky130_fd_sc_hd__inv_2 \inv[3039]/_0_  (.A(\inv_in[3039] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3040] ));
 sky130_fd_sc_hd__inv_2 \inv[303]/_0_  (.A(\inv_in[303] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[304] ));
 sky130_fd_sc_hd__inv_2 \inv[3040]/_0_  (.A(\inv_in[3040] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3041] ));
 sky130_fd_sc_hd__inv_2 \inv[3041]/_0_  (.A(\inv_in[3041] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3042] ));
 sky130_fd_sc_hd__inv_2 \inv[3042]/_0_  (.A(\inv_in[3042] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3043] ));
 sky130_fd_sc_hd__inv_2 \inv[3043]/_0_  (.A(\inv_in[3043] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3044] ));
 sky130_fd_sc_hd__inv_2 \inv[3044]/_0_  (.A(\inv_in[3044] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3045] ));
 sky130_fd_sc_hd__inv_2 \inv[3045]/_0_  (.A(\inv_in[3045] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3046] ));
 sky130_fd_sc_hd__inv_2 \inv[3046]/_0_  (.A(\inv_in[3046] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3047] ));
 sky130_fd_sc_hd__inv_2 \inv[3047]/_0_  (.A(\inv_in[3047] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3048] ));
 sky130_fd_sc_hd__inv_2 \inv[3048]/_0_  (.A(\inv_in[3048] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3049] ));
 sky130_fd_sc_hd__inv_2 \inv[3049]/_0_  (.A(\inv_in[3049] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3050] ));
 sky130_fd_sc_hd__inv_2 \inv[304]/_0_  (.A(\inv_in[304] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[305] ));
 sky130_fd_sc_hd__inv_2 \inv[3050]/_0_  (.A(\inv_in[3050] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3051] ));
 sky130_fd_sc_hd__inv_2 \inv[3051]/_0_  (.A(\inv_in[3051] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3052] ));
 sky130_fd_sc_hd__inv_2 \inv[3052]/_0_  (.A(\inv_in[3052] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3053] ));
 sky130_fd_sc_hd__inv_2 \inv[3053]/_0_  (.A(\inv_in[3053] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3054] ));
 sky130_fd_sc_hd__inv_2 \inv[3054]/_0_  (.A(\inv_in[3054] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3055] ));
 sky130_fd_sc_hd__inv_2 \inv[3055]/_0_  (.A(\inv_in[3055] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3056] ));
 sky130_fd_sc_hd__inv_2 \inv[3056]/_0_  (.A(\inv_in[3056] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3057] ));
 sky130_fd_sc_hd__inv_2 \inv[3057]/_0_  (.A(\inv_in[3057] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3058] ));
 sky130_fd_sc_hd__inv_2 \inv[3058]/_0_  (.A(\inv_in[3058] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3059] ));
 sky130_fd_sc_hd__inv_2 \inv[3059]/_0_  (.A(\inv_in[3059] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3060] ));
 sky130_fd_sc_hd__inv_2 \inv[305]/_0_  (.A(\inv_in[305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[306] ));
 sky130_fd_sc_hd__inv_2 \inv[3060]/_0_  (.A(\inv_in[3060] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3061] ));
 sky130_fd_sc_hd__inv_2 \inv[3061]/_0_  (.A(\inv_in[3061] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3062] ));
 sky130_fd_sc_hd__inv_2 \inv[3062]/_0_  (.A(\inv_in[3062] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3063] ));
 sky130_fd_sc_hd__inv_2 \inv[3063]/_0_  (.A(\inv_in[3063] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3064] ));
 sky130_fd_sc_hd__inv_2 \inv[3064]/_0_  (.A(\inv_in[3064] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3065] ));
 sky130_fd_sc_hd__inv_2 \inv[3065]/_0_  (.A(\inv_in[3065] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3066] ));
 sky130_fd_sc_hd__inv_2 \inv[3066]/_0_  (.A(\inv_in[3066] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3067] ));
 sky130_fd_sc_hd__inv_2 \inv[3067]/_0_  (.A(\inv_in[3067] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3068] ));
 sky130_fd_sc_hd__inv_2 \inv[3068]/_0_  (.A(\inv_in[3068] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3069] ));
 sky130_fd_sc_hd__inv_2 \inv[3069]/_0_  (.A(\inv_in[3069] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3070] ));
 sky130_fd_sc_hd__inv_2 \inv[306]/_0_  (.A(\inv_in[306] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[307] ));
 sky130_fd_sc_hd__inv_2 \inv[3070]/_0_  (.A(\inv_in[3070] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3071] ));
 sky130_fd_sc_hd__inv_2 \inv[3071]/_0_  (.A(\inv_in[3071] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3072] ));
 sky130_fd_sc_hd__inv_2 \inv[3072]/_0_  (.A(\inv_in[3072] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3073] ));
 sky130_fd_sc_hd__inv_2 \inv[3073]/_0_  (.A(\inv_in[3073] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3074] ));
 sky130_fd_sc_hd__inv_2 \inv[3074]/_0_  (.A(\inv_in[3074] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3075] ));
 sky130_fd_sc_hd__inv_2 \inv[3075]/_0_  (.A(\inv_in[3075] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3076] ));
 sky130_fd_sc_hd__inv_2 \inv[3076]/_0_  (.A(\inv_in[3076] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3077] ));
 sky130_fd_sc_hd__inv_2 \inv[3077]/_0_  (.A(\inv_in[3077] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3078] ));
 sky130_fd_sc_hd__inv_2 \inv[3078]/_0_  (.A(\inv_in[3078] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3079] ));
 sky130_fd_sc_hd__inv_2 \inv[3079]/_0_  (.A(\inv_in[3079] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3080] ));
 sky130_fd_sc_hd__inv_2 \inv[307]/_0_  (.A(\inv_in[307] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[308] ));
 sky130_fd_sc_hd__inv_2 \inv[3080]/_0_  (.A(\inv_in[3080] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3081] ));
 sky130_fd_sc_hd__inv_2 \inv[3081]/_0_  (.A(\inv_in[3081] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3082] ));
 sky130_fd_sc_hd__inv_2 \inv[3082]/_0_  (.A(\inv_in[3082] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3083] ));
 sky130_fd_sc_hd__inv_2 \inv[3083]/_0_  (.A(\inv_in[3083] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3084] ));
 sky130_fd_sc_hd__inv_2 \inv[3084]/_0_  (.A(\inv_in[3084] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3085] ));
 sky130_fd_sc_hd__inv_2 \inv[3085]/_0_  (.A(\inv_in[3085] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3086] ));
 sky130_fd_sc_hd__inv_2 \inv[3086]/_0_  (.A(\inv_in[3086] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3087] ));
 sky130_fd_sc_hd__inv_2 \inv[3087]/_0_  (.A(\inv_in[3087] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3088] ));
 sky130_fd_sc_hd__inv_2 \inv[3088]/_0_  (.A(\inv_in[3088] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3089] ));
 sky130_fd_sc_hd__inv_2 \inv[3089]/_0_  (.A(\inv_in[3089] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3090] ));
 sky130_fd_sc_hd__inv_2 \inv[308]/_0_  (.A(\inv_in[308] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[309] ));
 sky130_fd_sc_hd__inv_2 \inv[3090]/_0_  (.A(\inv_in[3090] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3091] ));
 sky130_fd_sc_hd__inv_2 \inv[3091]/_0_  (.A(\inv_in[3091] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3092] ));
 sky130_fd_sc_hd__inv_2 \inv[3092]/_0_  (.A(\inv_in[3092] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3093] ));
 sky130_fd_sc_hd__inv_2 \inv[3093]/_0_  (.A(\inv_in[3093] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3094] ));
 sky130_fd_sc_hd__inv_2 \inv[3094]/_0_  (.A(\inv_in[3094] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3095] ));
 sky130_fd_sc_hd__inv_2 \inv[3095]/_0_  (.A(\inv_in[3095] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3096] ));
 sky130_fd_sc_hd__inv_2 \inv[3096]/_0_  (.A(\inv_in[3096] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3097] ));
 sky130_fd_sc_hd__inv_2 \inv[3097]/_0_  (.A(\inv_in[3097] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3098] ));
 sky130_fd_sc_hd__inv_2 \inv[3098]/_0_  (.A(\inv_in[3098] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3099] ));
 sky130_fd_sc_hd__inv_2 \inv[3099]/_0_  (.A(\inv_in[3099] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3100] ));
 sky130_fd_sc_hd__inv_2 \inv[309]/_0_  (.A(\inv_in[309] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[310] ));
 sky130_fd_sc_hd__inv_2 \inv[30]/_0_  (.A(\inv_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[31] ));
 sky130_fd_sc_hd__inv_2 \inv[3100]/_0_  (.A(\inv_in[3100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3101] ));
 sky130_fd_sc_hd__inv_2 \inv[3101]/_0_  (.A(\inv_in[3101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3102] ));
 sky130_fd_sc_hd__inv_2 \inv[3102]/_0_  (.A(\inv_in[3102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3103] ));
 sky130_fd_sc_hd__inv_2 \inv[3103]/_0_  (.A(\inv_in[3103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3104] ));
 sky130_fd_sc_hd__inv_2 \inv[3104]/_0_  (.A(\inv_in[3104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3105] ));
 sky130_fd_sc_hd__inv_2 \inv[3105]/_0_  (.A(\inv_in[3105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3106] ));
 sky130_fd_sc_hd__inv_2 \inv[3106]/_0_  (.A(\inv_in[3106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3107] ));
 sky130_fd_sc_hd__inv_2 \inv[3107]/_0_  (.A(\inv_in[3107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3108] ));
 sky130_fd_sc_hd__inv_2 \inv[3108]/_0_  (.A(\inv_in[3108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3109] ));
 sky130_fd_sc_hd__inv_2 \inv[3109]/_0_  (.A(\inv_in[3109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3110] ));
 sky130_fd_sc_hd__inv_2 \inv[310]/_0_  (.A(\inv_in[310] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[311] ));
 sky130_fd_sc_hd__inv_2 \inv[3110]/_0_  (.A(\inv_in[3110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3111] ));
 sky130_fd_sc_hd__inv_2 \inv[3111]/_0_  (.A(\inv_in[3111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3112] ));
 sky130_fd_sc_hd__inv_2 \inv[3112]/_0_  (.A(\inv_in[3112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3113] ));
 sky130_fd_sc_hd__inv_2 \inv[3113]/_0_  (.A(\inv_in[3113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3114] ));
 sky130_fd_sc_hd__inv_2 \inv[3114]/_0_  (.A(\inv_in[3114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3115] ));
 sky130_fd_sc_hd__inv_2 \inv[3115]/_0_  (.A(\inv_in[3115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3116] ));
 sky130_fd_sc_hd__inv_2 \inv[3116]/_0_  (.A(\inv_in[3116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3117] ));
 sky130_fd_sc_hd__inv_2 \inv[3117]/_0_  (.A(\inv_in[3117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3118] ));
 sky130_fd_sc_hd__inv_2 \inv[3118]/_0_  (.A(\inv_in[3118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3119] ));
 sky130_fd_sc_hd__inv_2 \inv[3119]/_0_  (.A(\inv_in[3119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3120] ));
 sky130_fd_sc_hd__inv_2 \inv[311]/_0_  (.A(\inv_in[311] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[312] ));
 sky130_fd_sc_hd__inv_2 \inv[3120]/_0_  (.A(\inv_in[3120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3121] ));
 sky130_fd_sc_hd__inv_2 \inv[3121]/_0_  (.A(\inv_in[3121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3122] ));
 sky130_fd_sc_hd__inv_2 \inv[3122]/_0_  (.A(\inv_in[3122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3123] ));
 sky130_fd_sc_hd__inv_2 \inv[3123]/_0_  (.A(\inv_in[3123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3124] ));
 sky130_fd_sc_hd__inv_2 \inv[3124]/_0_  (.A(\inv_in[3124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3125] ));
 sky130_fd_sc_hd__inv_2 \inv[3125]/_0_  (.A(\inv_in[3125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3126] ));
 sky130_fd_sc_hd__inv_2 \inv[3126]/_0_  (.A(\inv_in[3126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3127] ));
 sky130_fd_sc_hd__inv_2 \inv[3127]/_0_  (.A(\inv_in[3127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3128] ));
 sky130_fd_sc_hd__inv_2 \inv[3128]/_0_  (.A(\inv_in[3128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3129] ));
 sky130_fd_sc_hd__inv_2 \inv[3129]/_0_  (.A(\inv_in[3129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3130] ));
 sky130_fd_sc_hd__inv_2 \inv[312]/_0_  (.A(\inv_in[312] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[313] ));
 sky130_fd_sc_hd__inv_2 \inv[3130]/_0_  (.A(\inv_in[3130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3131] ));
 sky130_fd_sc_hd__inv_2 \inv[3131]/_0_  (.A(\inv_in[3131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3132] ));
 sky130_fd_sc_hd__inv_2 \inv[3132]/_0_  (.A(\inv_in[3132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3133] ));
 sky130_fd_sc_hd__inv_2 \inv[3133]/_0_  (.A(\inv_in[3133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3134] ));
 sky130_fd_sc_hd__inv_2 \inv[3134]/_0_  (.A(\inv_in[3134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3135] ));
 sky130_fd_sc_hd__inv_2 \inv[3135]/_0_  (.A(\inv_in[3135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3136] ));
 sky130_fd_sc_hd__inv_2 \inv[3136]/_0_  (.A(\inv_in[3136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3137] ));
 sky130_fd_sc_hd__inv_2 \inv[3137]/_0_  (.A(\inv_in[3137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3138] ));
 sky130_fd_sc_hd__inv_2 \inv[3138]/_0_  (.A(\inv_in[3138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3139] ));
 sky130_fd_sc_hd__inv_2 \inv[3139]/_0_  (.A(\inv_in[3139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3140] ));
 sky130_fd_sc_hd__inv_2 \inv[313]/_0_  (.A(\inv_in[313] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[314] ));
 sky130_fd_sc_hd__inv_2 \inv[3140]/_0_  (.A(\inv_in[3140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3141] ));
 sky130_fd_sc_hd__inv_2 \inv[3141]/_0_  (.A(\inv_in[3141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3142] ));
 sky130_fd_sc_hd__inv_2 \inv[3142]/_0_  (.A(\inv_in[3142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3143] ));
 sky130_fd_sc_hd__inv_2 \inv[3143]/_0_  (.A(\inv_in[3143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3144] ));
 sky130_fd_sc_hd__inv_2 \inv[3144]/_0_  (.A(\inv_in[3144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3145] ));
 sky130_fd_sc_hd__inv_2 \inv[3145]/_0_  (.A(\inv_in[3145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3146] ));
 sky130_fd_sc_hd__inv_2 \inv[3146]/_0_  (.A(\inv_in[3146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3147] ));
 sky130_fd_sc_hd__inv_2 \inv[3147]/_0_  (.A(\inv_in[3147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3148] ));
 sky130_fd_sc_hd__inv_2 \inv[3148]/_0_  (.A(\inv_in[3148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3149] ));
 sky130_fd_sc_hd__inv_2 \inv[3149]/_0_  (.A(\inv_in[3149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3150] ));
 sky130_fd_sc_hd__inv_2 \inv[314]/_0_  (.A(\inv_in[314] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[315] ));
 sky130_fd_sc_hd__inv_2 \inv[3150]/_0_  (.A(\inv_in[3150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3151] ));
 sky130_fd_sc_hd__inv_2 \inv[3151]/_0_  (.A(\inv_in[3151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3152] ));
 sky130_fd_sc_hd__inv_2 \inv[3152]/_0_  (.A(\inv_in[3152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3153] ));
 sky130_fd_sc_hd__inv_2 \inv[3153]/_0_  (.A(\inv_in[3153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3154] ));
 sky130_fd_sc_hd__inv_2 \inv[3154]/_0_  (.A(\inv_in[3154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3155] ));
 sky130_fd_sc_hd__inv_2 \inv[3155]/_0_  (.A(\inv_in[3155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3156] ));
 sky130_fd_sc_hd__inv_2 \inv[3156]/_0_  (.A(\inv_in[3156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3157] ));
 sky130_fd_sc_hd__inv_2 \inv[3157]/_0_  (.A(\inv_in[3157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3158] ));
 sky130_fd_sc_hd__inv_2 \inv[3158]/_0_  (.A(\inv_in[3158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3159] ));
 sky130_fd_sc_hd__inv_2 \inv[3159]/_0_  (.A(\inv_in[3159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3160] ));
 sky130_fd_sc_hd__inv_2 \inv[315]/_0_  (.A(\inv_in[315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[316] ));
 sky130_fd_sc_hd__inv_2 \inv[3160]/_0_  (.A(\inv_in[3160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3161] ));
 sky130_fd_sc_hd__inv_2 \inv[3161]/_0_  (.A(\inv_in[3161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3162] ));
 sky130_fd_sc_hd__inv_2 \inv[3162]/_0_  (.A(\inv_in[3162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3163] ));
 sky130_fd_sc_hd__inv_2 \inv[3163]/_0_  (.A(\inv_in[3163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3164] ));
 sky130_fd_sc_hd__inv_2 \inv[3164]/_0_  (.A(\inv_in[3164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3165] ));
 sky130_fd_sc_hd__inv_2 \inv[3165]/_0_  (.A(\inv_in[3165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3166] ));
 sky130_fd_sc_hd__inv_2 \inv[3166]/_0_  (.A(\inv_in[3166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3167] ));
 sky130_fd_sc_hd__inv_2 \inv[3167]/_0_  (.A(\inv_in[3167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3168] ));
 sky130_fd_sc_hd__inv_2 \inv[3168]/_0_  (.A(\inv_in[3168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3169] ));
 sky130_fd_sc_hd__inv_2 \inv[3169]/_0_  (.A(\inv_in[3169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3170] ));
 sky130_fd_sc_hd__inv_2 \inv[316]/_0_  (.A(\inv_in[316] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[317] ));
 sky130_fd_sc_hd__inv_2 \inv[3170]/_0_  (.A(\inv_in[3170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3171] ));
 sky130_fd_sc_hd__inv_2 \inv[3171]/_0_  (.A(\inv_in[3171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3172] ));
 sky130_fd_sc_hd__inv_2 \inv[3172]/_0_  (.A(\inv_in[3172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3173] ));
 sky130_fd_sc_hd__inv_2 \inv[3173]/_0_  (.A(\inv_in[3173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3174] ));
 sky130_fd_sc_hd__inv_2 \inv[3174]/_0_  (.A(\inv_in[3174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3175] ));
 sky130_fd_sc_hd__inv_2 \inv[3175]/_0_  (.A(\inv_in[3175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3176] ));
 sky130_fd_sc_hd__inv_2 \inv[3176]/_0_  (.A(\inv_in[3176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3177] ));
 sky130_fd_sc_hd__inv_2 \inv[3177]/_0_  (.A(\inv_in[3177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3178] ));
 sky130_fd_sc_hd__inv_2 \inv[3178]/_0_  (.A(\inv_in[3178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3179] ));
 sky130_fd_sc_hd__inv_2 \inv[3179]/_0_  (.A(\inv_in[3179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3180] ));
 sky130_fd_sc_hd__inv_2 \inv[317]/_0_  (.A(\inv_in[317] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[318] ));
 sky130_fd_sc_hd__inv_2 \inv[3180]/_0_  (.A(\inv_in[3180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3181] ));
 sky130_fd_sc_hd__inv_2 \inv[3181]/_0_  (.A(\inv_in[3181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3182] ));
 sky130_fd_sc_hd__inv_2 \inv[3182]/_0_  (.A(\inv_in[3182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3183] ));
 sky130_fd_sc_hd__inv_2 \inv[3183]/_0_  (.A(\inv_in[3183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3184] ));
 sky130_fd_sc_hd__inv_2 \inv[3184]/_0_  (.A(\inv_in[3184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3185] ));
 sky130_fd_sc_hd__inv_2 \inv[3185]/_0_  (.A(\inv_in[3185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3186] ));
 sky130_fd_sc_hd__inv_2 \inv[3186]/_0_  (.A(\inv_in[3186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3187] ));
 sky130_fd_sc_hd__inv_2 \inv[3187]/_0_  (.A(\inv_in[3187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3188] ));
 sky130_fd_sc_hd__inv_2 \inv[3188]/_0_  (.A(\inv_in[3188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3189] ));
 sky130_fd_sc_hd__inv_2 \inv[3189]/_0_  (.A(\inv_in[3189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3190] ));
 sky130_fd_sc_hd__inv_2 \inv[318]/_0_  (.A(\inv_in[318] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[319] ));
 sky130_fd_sc_hd__inv_2 \inv[3190]/_0_  (.A(\inv_in[3190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3191] ));
 sky130_fd_sc_hd__inv_2 \inv[3191]/_0_  (.A(\inv_in[3191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3192] ));
 sky130_fd_sc_hd__inv_2 \inv[3192]/_0_  (.A(\inv_in[3192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3193] ));
 sky130_fd_sc_hd__inv_2 \inv[3193]/_0_  (.A(\inv_in[3193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3194] ));
 sky130_fd_sc_hd__inv_2 \inv[3194]/_0_  (.A(\inv_in[3194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3195] ));
 sky130_fd_sc_hd__inv_2 \inv[3195]/_0_  (.A(\inv_in[3195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3196] ));
 sky130_fd_sc_hd__inv_2 \inv[3196]/_0_  (.A(\inv_in[3196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3197] ));
 sky130_fd_sc_hd__inv_2 \inv[3197]/_0_  (.A(\inv_in[3197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3198] ));
 sky130_fd_sc_hd__inv_2 \inv[3198]/_0_  (.A(\inv_in[3198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3199] ));
 sky130_fd_sc_hd__inv_2 \inv[3199]/_0_  (.A(\inv_in[3199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3200] ));
 sky130_fd_sc_hd__inv_2 \inv[319]/_0_  (.A(\inv_in[319] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[320] ));
 sky130_fd_sc_hd__inv_2 \inv[31]/_0_  (.A(\inv_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[32] ));
 sky130_fd_sc_hd__inv_2 \inv[3200]/_0_  (.A(\inv_in[3200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3201] ));
 sky130_fd_sc_hd__inv_2 \inv[3201]/_0_  (.A(\inv_in[3201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3202] ));
 sky130_fd_sc_hd__inv_2 \inv[3202]/_0_  (.A(\inv_in[3202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3203] ));
 sky130_fd_sc_hd__inv_2 \inv[3203]/_0_  (.A(\inv_in[3203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3204] ));
 sky130_fd_sc_hd__inv_2 \inv[3204]/_0_  (.A(\inv_in[3204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3205] ));
 sky130_fd_sc_hd__inv_2 \inv[3205]/_0_  (.A(\inv_in[3205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3206] ));
 sky130_fd_sc_hd__inv_2 \inv[3206]/_0_  (.A(\inv_in[3206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3207] ));
 sky130_fd_sc_hd__inv_2 \inv[3207]/_0_  (.A(\inv_in[3207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3208] ));
 sky130_fd_sc_hd__inv_2 \inv[3208]/_0_  (.A(\inv_in[3208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3209] ));
 sky130_fd_sc_hd__inv_2 \inv[3209]/_0_  (.A(\inv_in[3209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3210] ));
 sky130_fd_sc_hd__inv_2 \inv[320]/_0_  (.A(\inv_in[320] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[321] ));
 sky130_fd_sc_hd__inv_2 \inv[3210]/_0_  (.A(\inv_in[3210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3211] ));
 sky130_fd_sc_hd__inv_2 \inv[3211]/_0_  (.A(\inv_in[3211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3212] ));
 sky130_fd_sc_hd__inv_2 \inv[3212]/_0_  (.A(\inv_in[3212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3213] ));
 sky130_fd_sc_hd__inv_2 \inv[3213]/_0_  (.A(\inv_in[3213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3214] ));
 sky130_fd_sc_hd__inv_2 \inv[3214]/_0_  (.A(\inv_in[3214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3215] ));
 sky130_fd_sc_hd__inv_2 \inv[3215]/_0_  (.A(\inv_in[3215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3216] ));
 sky130_fd_sc_hd__inv_2 \inv[3216]/_0_  (.A(\inv_in[3216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3217] ));
 sky130_fd_sc_hd__inv_2 \inv[3217]/_0_  (.A(\inv_in[3217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3218] ));
 sky130_fd_sc_hd__inv_2 \inv[3218]/_0_  (.A(\inv_in[3218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3219] ));
 sky130_fd_sc_hd__inv_2 \inv[3219]/_0_  (.A(\inv_in[3219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3220] ));
 sky130_fd_sc_hd__inv_2 \inv[321]/_0_  (.A(\inv_in[321] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[322] ));
 sky130_fd_sc_hd__inv_2 \inv[3220]/_0_  (.A(\inv_in[3220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3221] ));
 sky130_fd_sc_hd__inv_2 \inv[3221]/_0_  (.A(\inv_in[3221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3222] ));
 sky130_fd_sc_hd__inv_2 \inv[3222]/_0_  (.A(\inv_in[3222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3223] ));
 sky130_fd_sc_hd__inv_2 \inv[3223]/_0_  (.A(\inv_in[3223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3224] ));
 sky130_fd_sc_hd__inv_2 \inv[3224]/_0_  (.A(\inv_in[3224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3225] ));
 sky130_fd_sc_hd__inv_2 \inv[3225]/_0_  (.A(\inv_in[3225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3226] ));
 sky130_fd_sc_hd__inv_2 \inv[3226]/_0_  (.A(\inv_in[3226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3227] ));
 sky130_fd_sc_hd__inv_2 \inv[3227]/_0_  (.A(\inv_in[3227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3228] ));
 sky130_fd_sc_hd__inv_2 \inv[3228]/_0_  (.A(\inv_in[3228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3229] ));
 sky130_fd_sc_hd__inv_2 \inv[3229]/_0_  (.A(\inv_in[3229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3230] ));
 sky130_fd_sc_hd__inv_2 \inv[322]/_0_  (.A(\inv_in[322] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[323] ));
 sky130_fd_sc_hd__inv_2 \inv[3230]/_0_  (.A(\inv_in[3230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3231] ));
 sky130_fd_sc_hd__inv_2 \inv[3231]/_0_  (.A(\inv_in[3231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3232] ));
 sky130_fd_sc_hd__inv_2 \inv[3232]/_0_  (.A(\inv_in[3232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3233] ));
 sky130_fd_sc_hd__inv_2 \inv[3233]/_0_  (.A(\inv_in[3233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3234] ));
 sky130_fd_sc_hd__inv_2 \inv[3234]/_0_  (.A(\inv_in[3234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3235] ));
 sky130_fd_sc_hd__inv_2 \inv[3235]/_0_  (.A(\inv_in[3235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3236] ));
 sky130_fd_sc_hd__inv_2 \inv[3236]/_0_  (.A(\inv_in[3236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3237] ));
 sky130_fd_sc_hd__inv_2 \inv[3237]/_0_  (.A(\inv_in[3237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3238] ));
 sky130_fd_sc_hd__inv_2 \inv[3238]/_0_  (.A(\inv_in[3238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3239] ));
 sky130_fd_sc_hd__inv_2 \inv[3239]/_0_  (.A(\inv_in[3239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3240] ));
 sky130_fd_sc_hd__inv_2 \inv[323]/_0_  (.A(\inv_in[323] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[324] ));
 sky130_fd_sc_hd__inv_2 \inv[3240]/_0_  (.A(\inv_in[3240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3241] ));
 sky130_fd_sc_hd__inv_2 \inv[3241]/_0_  (.A(\inv_in[3241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3242] ));
 sky130_fd_sc_hd__inv_2 \inv[3242]/_0_  (.A(\inv_in[3242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3243] ));
 sky130_fd_sc_hd__inv_2 \inv[3243]/_0_  (.A(\inv_in[3243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3244] ));
 sky130_fd_sc_hd__inv_2 \inv[3244]/_0_  (.A(\inv_in[3244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3245] ));
 sky130_fd_sc_hd__inv_2 \inv[3245]/_0_  (.A(\inv_in[3245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3246] ));
 sky130_fd_sc_hd__inv_2 \inv[3246]/_0_  (.A(\inv_in[3246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3247] ));
 sky130_fd_sc_hd__inv_2 \inv[3247]/_0_  (.A(\inv_in[3247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3248] ));
 sky130_fd_sc_hd__inv_2 \inv[3248]/_0_  (.A(\inv_in[3248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3249] ));
 sky130_fd_sc_hd__inv_2 \inv[3249]/_0_  (.A(\inv_in[3249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3250] ));
 sky130_fd_sc_hd__inv_2 \inv[324]/_0_  (.A(\inv_in[324] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[325] ));
 sky130_fd_sc_hd__inv_2 \inv[3250]/_0_  (.A(\inv_in[3250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3251] ));
 sky130_fd_sc_hd__inv_2 \inv[3251]/_0_  (.A(\inv_in[3251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3252] ));
 sky130_fd_sc_hd__inv_2 \inv[3252]/_0_  (.A(\inv_in[3252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3253] ));
 sky130_fd_sc_hd__inv_2 \inv[3253]/_0_  (.A(\inv_in[3253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3254] ));
 sky130_fd_sc_hd__inv_2 \inv[3254]/_0_  (.A(\inv_in[3254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3255] ));
 sky130_fd_sc_hd__inv_2 \inv[3255]/_0_  (.A(\inv_in[3255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3256] ));
 sky130_fd_sc_hd__inv_2 \inv[3256]/_0_  (.A(\inv_in[3256] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3257] ));
 sky130_fd_sc_hd__inv_2 \inv[3257]/_0_  (.A(\inv_in[3257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3258] ));
 sky130_fd_sc_hd__inv_2 \inv[3258]/_0_  (.A(\inv_in[3258] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3259] ));
 sky130_fd_sc_hd__inv_2 \inv[3259]/_0_  (.A(\inv_in[3259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3260] ));
 sky130_fd_sc_hd__inv_2 \inv[325]/_0_  (.A(\inv_in[325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[326] ));
 sky130_fd_sc_hd__inv_2 \inv[3260]/_0_  (.A(\inv_in[3260] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3261] ));
 sky130_fd_sc_hd__inv_2 \inv[3261]/_0_  (.A(\inv_in[3261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3262] ));
 sky130_fd_sc_hd__inv_2 \inv[3262]/_0_  (.A(\inv_in[3262] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3263] ));
 sky130_fd_sc_hd__inv_2 \inv[3263]/_0_  (.A(\inv_in[3263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3264] ));
 sky130_fd_sc_hd__inv_2 \inv[3264]/_0_  (.A(\inv_in[3264] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3265] ));
 sky130_fd_sc_hd__inv_2 \inv[3265]/_0_  (.A(\inv_in[3265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3266] ));
 sky130_fd_sc_hd__inv_2 \inv[3266]/_0_  (.A(\inv_in[3266] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3267] ));
 sky130_fd_sc_hd__inv_2 \inv[3267]/_0_  (.A(\inv_in[3267] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3268] ));
 sky130_fd_sc_hd__inv_2 \inv[3268]/_0_  (.A(\inv_in[3268] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3269] ));
 sky130_fd_sc_hd__inv_2 \inv[3269]/_0_  (.A(\inv_in[3269] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3270] ));
 sky130_fd_sc_hd__inv_2 \inv[326]/_0_  (.A(\inv_in[326] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[327] ));
 sky130_fd_sc_hd__inv_2 \inv[3270]/_0_  (.A(\inv_in[3270] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3271] ));
 sky130_fd_sc_hd__inv_2 \inv[3271]/_0_  (.A(\inv_in[3271] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3272] ));
 sky130_fd_sc_hd__inv_2 \inv[3272]/_0_  (.A(\inv_in[3272] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3273] ));
 sky130_fd_sc_hd__inv_2 \inv[3273]/_0_  (.A(\inv_in[3273] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3274] ));
 sky130_fd_sc_hd__inv_2 \inv[3274]/_0_  (.A(\inv_in[3274] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3275] ));
 sky130_fd_sc_hd__inv_2 \inv[3275]/_0_  (.A(\inv_in[3275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3276] ));
 sky130_fd_sc_hd__inv_2 \inv[3276]/_0_  (.A(\inv_in[3276] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3277] ));
 sky130_fd_sc_hd__inv_2 \inv[3277]/_0_  (.A(\inv_in[3277] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3278] ));
 sky130_fd_sc_hd__inv_2 \inv[3278]/_0_  (.A(\inv_in[3278] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3279] ));
 sky130_fd_sc_hd__inv_2 \inv[3279]/_0_  (.A(\inv_in[3279] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3280] ));
 sky130_fd_sc_hd__inv_2 \inv[327]/_0_  (.A(\inv_in[327] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[328] ));
 sky130_fd_sc_hd__inv_2 \inv[3280]/_0_  (.A(\inv_in[3280] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3281] ));
 sky130_fd_sc_hd__inv_2 \inv[3281]/_0_  (.A(\inv_in[3281] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3282] ));
 sky130_fd_sc_hd__inv_2 \inv[3282]/_0_  (.A(\inv_in[3282] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3283] ));
 sky130_fd_sc_hd__inv_2 \inv[3283]/_0_  (.A(\inv_in[3283] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3284] ));
 sky130_fd_sc_hd__inv_2 \inv[3284]/_0_  (.A(\inv_in[3284] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3285] ));
 sky130_fd_sc_hd__inv_2 \inv[3285]/_0_  (.A(\inv_in[3285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3286] ));
 sky130_fd_sc_hd__inv_2 \inv[3286]/_0_  (.A(\inv_in[3286] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3287] ));
 sky130_fd_sc_hd__inv_2 \inv[3287]/_0_  (.A(\inv_in[3287] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3288] ));
 sky130_fd_sc_hd__inv_2 \inv[3288]/_0_  (.A(\inv_in[3288] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3289] ));
 sky130_fd_sc_hd__inv_2 \inv[3289]/_0_  (.A(\inv_in[3289] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3290] ));
 sky130_fd_sc_hd__inv_2 \inv[328]/_0_  (.A(\inv_in[328] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[329] ));
 sky130_fd_sc_hd__inv_2 \inv[3290]/_0_  (.A(\inv_in[3290] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3291] ));
 sky130_fd_sc_hd__inv_2 \inv[3291]/_0_  (.A(\inv_in[3291] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3292] ));
 sky130_fd_sc_hd__inv_2 \inv[3292]/_0_  (.A(\inv_in[3292] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3293] ));
 sky130_fd_sc_hd__inv_2 \inv[3293]/_0_  (.A(\inv_in[3293] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3294] ));
 sky130_fd_sc_hd__inv_2 \inv[3294]/_0_  (.A(\inv_in[3294] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3295] ));
 sky130_fd_sc_hd__inv_2 \inv[3295]/_0_  (.A(\inv_in[3295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3296] ));
 sky130_fd_sc_hd__inv_2 \inv[3296]/_0_  (.A(\inv_in[3296] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3297] ));
 sky130_fd_sc_hd__inv_2 \inv[3297]/_0_  (.A(\inv_in[3297] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3298] ));
 sky130_fd_sc_hd__inv_2 \inv[3298]/_0_  (.A(\inv_in[3298] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3299] ));
 sky130_fd_sc_hd__inv_2 \inv[3299]/_0_  (.A(\inv_in[3299] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3300] ));
 sky130_fd_sc_hd__inv_2 \inv[329]/_0_  (.A(\inv_in[329] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[330] ));
 sky130_fd_sc_hd__inv_2 \inv[32]/_0_  (.A(\inv_in[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[33] ));
 sky130_fd_sc_hd__inv_2 \inv[3300]/_0_  (.A(\inv_in[3300] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3301] ));
 sky130_fd_sc_hd__inv_2 \inv[3301]/_0_  (.A(\inv_in[3301] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3302] ));
 sky130_fd_sc_hd__inv_2 \inv[3302]/_0_  (.A(\inv_in[3302] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3303] ));
 sky130_fd_sc_hd__inv_2 \inv[3303]/_0_  (.A(\inv_in[3303] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3304] ));
 sky130_fd_sc_hd__inv_2 \inv[3304]/_0_  (.A(\inv_in[3304] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3305] ));
 sky130_fd_sc_hd__inv_2 \inv[3305]/_0_  (.A(\inv_in[3305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3306] ));
 sky130_fd_sc_hd__inv_2 \inv[3306]/_0_  (.A(\inv_in[3306] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3307] ));
 sky130_fd_sc_hd__inv_2 \inv[3307]/_0_  (.A(\inv_in[3307] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3308] ));
 sky130_fd_sc_hd__inv_2 \inv[3308]/_0_  (.A(\inv_in[3308] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3309] ));
 sky130_fd_sc_hd__inv_2 \inv[3309]/_0_  (.A(\inv_in[3309] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3310] ));
 sky130_fd_sc_hd__inv_2 \inv[330]/_0_  (.A(\inv_in[330] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[331] ));
 sky130_fd_sc_hd__inv_2 \inv[3310]/_0_  (.A(\inv_in[3310] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3311] ));
 sky130_fd_sc_hd__inv_2 \inv[3311]/_0_  (.A(\inv_in[3311] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3312] ));
 sky130_fd_sc_hd__inv_2 \inv[3312]/_0_  (.A(\inv_in[3312] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3313] ));
 sky130_fd_sc_hd__inv_2 \inv[3313]/_0_  (.A(\inv_in[3313] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3314] ));
 sky130_fd_sc_hd__inv_2 \inv[3314]/_0_  (.A(\inv_in[3314] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3315] ));
 sky130_fd_sc_hd__inv_2 \inv[3315]/_0_  (.A(\inv_in[3315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3316] ));
 sky130_fd_sc_hd__inv_2 \inv[3316]/_0_  (.A(\inv_in[3316] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3317] ));
 sky130_fd_sc_hd__inv_2 \inv[3317]/_0_  (.A(\inv_in[3317] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3318] ));
 sky130_fd_sc_hd__inv_2 \inv[3318]/_0_  (.A(\inv_in[3318] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3319] ));
 sky130_fd_sc_hd__inv_2 \inv[3319]/_0_  (.A(\inv_in[3319] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3320] ));
 sky130_fd_sc_hd__inv_2 \inv[331]/_0_  (.A(\inv_in[331] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[332] ));
 sky130_fd_sc_hd__inv_2 \inv[3320]/_0_  (.A(\inv_in[3320] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3321] ));
 sky130_fd_sc_hd__inv_2 \inv[3321]/_0_  (.A(\inv_in[3321] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3322] ));
 sky130_fd_sc_hd__inv_2 \inv[3322]/_0_  (.A(\inv_in[3322] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3323] ));
 sky130_fd_sc_hd__inv_2 \inv[3323]/_0_  (.A(\inv_in[3323] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3324] ));
 sky130_fd_sc_hd__inv_2 \inv[3324]/_0_  (.A(\inv_in[3324] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3325] ));
 sky130_fd_sc_hd__inv_2 \inv[3325]/_0_  (.A(\inv_in[3325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3326] ));
 sky130_fd_sc_hd__inv_2 \inv[3326]/_0_  (.A(\inv_in[3326] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3327] ));
 sky130_fd_sc_hd__inv_2 \inv[3327]/_0_  (.A(\inv_in[3327] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3328] ));
 sky130_fd_sc_hd__inv_2 \inv[3328]/_0_  (.A(\inv_in[3328] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3329] ));
 sky130_fd_sc_hd__inv_2 \inv[3329]/_0_  (.A(\inv_in[3329] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3330] ));
 sky130_fd_sc_hd__inv_2 \inv[332]/_0_  (.A(\inv_in[332] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[333] ));
 sky130_fd_sc_hd__inv_2 \inv[3330]/_0_  (.A(\inv_in[3330] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3331] ));
 sky130_fd_sc_hd__inv_2 \inv[3331]/_0_  (.A(\inv_in[3331] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3332] ));
 sky130_fd_sc_hd__inv_2 \inv[3332]/_0_  (.A(\inv_in[3332] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3333] ));
 sky130_fd_sc_hd__inv_2 \inv[3333]/_0_  (.A(\inv_in[3333] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3334] ));
 sky130_fd_sc_hd__inv_2 \inv[3334]/_0_  (.A(\inv_in[3334] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3335] ));
 sky130_fd_sc_hd__inv_2 \inv[3335]/_0_  (.A(\inv_in[3335] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3336] ));
 sky130_fd_sc_hd__inv_2 \inv[3336]/_0_  (.A(\inv_in[3336] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3337] ));
 sky130_fd_sc_hd__inv_2 \inv[3337]/_0_  (.A(\inv_in[3337] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3338] ));
 sky130_fd_sc_hd__inv_2 \inv[3338]/_0_  (.A(\inv_in[3338] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3339] ));
 sky130_fd_sc_hd__inv_2 \inv[3339]/_0_  (.A(\inv_in[3339] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3340] ));
 sky130_fd_sc_hd__inv_2 \inv[333]/_0_  (.A(\inv_in[333] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[334] ));
 sky130_fd_sc_hd__inv_2 \inv[3340]/_0_  (.A(\inv_in[3340] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3341] ));
 sky130_fd_sc_hd__inv_2 \inv[3341]/_0_  (.A(\inv_in[3341] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3342] ));
 sky130_fd_sc_hd__inv_2 \inv[3342]/_0_  (.A(\inv_in[3342] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3343] ));
 sky130_fd_sc_hd__inv_2 \inv[3343]/_0_  (.A(\inv_in[3343] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3344] ));
 sky130_fd_sc_hd__inv_2 \inv[3344]/_0_  (.A(\inv_in[3344] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3345] ));
 sky130_fd_sc_hd__inv_2 \inv[3345]/_0_  (.A(\inv_in[3345] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3346] ));
 sky130_fd_sc_hd__inv_2 \inv[3346]/_0_  (.A(\inv_in[3346] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3347] ));
 sky130_fd_sc_hd__inv_2 \inv[3347]/_0_  (.A(\inv_in[3347] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3348] ));
 sky130_fd_sc_hd__inv_2 \inv[3348]/_0_  (.A(\inv_in[3348] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3349] ));
 sky130_fd_sc_hd__inv_2 \inv[3349]/_0_  (.A(\inv_in[3349] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3350] ));
 sky130_fd_sc_hd__inv_2 \inv[334]/_0_  (.A(\inv_in[334] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[335] ));
 sky130_fd_sc_hd__inv_2 \inv[3350]/_0_  (.A(\inv_in[3350] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3351] ));
 sky130_fd_sc_hd__inv_2 \inv[3351]/_0_  (.A(\inv_in[3351] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3352] ));
 sky130_fd_sc_hd__inv_2 \inv[3352]/_0_  (.A(\inv_in[3352] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3353] ));
 sky130_fd_sc_hd__inv_2 \inv[3353]/_0_  (.A(\inv_in[3353] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3354] ));
 sky130_fd_sc_hd__inv_2 \inv[3354]/_0_  (.A(\inv_in[3354] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3355] ));
 sky130_fd_sc_hd__inv_2 \inv[3355]/_0_  (.A(\inv_in[3355] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3356] ));
 sky130_fd_sc_hd__inv_2 \inv[3356]/_0_  (.A(\inv_in[3356] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3357] ));
 sky130_fd_sc_hd__inv_2 \inv[3357]/_0_  (.A(\inv_in[3357] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3358] ));
 sky130_fd_sc_hd__inv_2 \inv[3358]/_0_  (.A(\inv_in[3358] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3359] ));
 sky130_fd_sc_hd__inv_2 \inv[3359]/_0_  (.A(\inv_in[3359] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3360] ));
 sky130_fd_sc_hd__inv_2 \inv[335]/_0_  (.A(\inv_in[335] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[336] ));
 sky130_fd_sc_hd__inv_2 \inv[3360]/_0_  (.A(\inv_in[3360] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3361] ));
 sky130_fd_sc_hd__inv_2 \inv[3361]/_0_  (.A(\inv_in[3361] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3362] ));
 sky130_fd_sc_hd__inv_2 \inv[3362]/_0_  (.A(\inv_in[3362] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3363] ));
 sky130_fd_sc_hd__inv_2 \inv[3363]/_0_  (.A(\inv_in[3363] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3364] ));
 sky130_fd_sc_hd__inv_2 \inv[3364]/_0_  (.A(\inv_in[3364] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3365] ));
 sky130_fd_sc_hd__inv_2 \inv[3365]/_0_  (.A(\inv_in[3365] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3366] ));
 sky130_fd_sc_hd__inv_2 \inv[3366]/_0_  (.A(\inv_in[3366] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3367] ));
 sky130_fd_sc_hd__inv_2 \inv[3367]/_0_  (.A(\inv_in[3367] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3368] ));
 sky130_fd_sc_hd__inv_2 \inv[3368]/_0_  (.A(\inv_in[3368] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3369] ));
 sky130_fd_sc_hd__inv_2 \inv[3369]/_0_  (.A(\inv_in[3369] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3370] ));
 sky130_fd_sc_hd__inv_2 \inv[336]/_0_  (.A(\inv_in[336] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[337] ));
 sky130_fd_sc_hd__inv_2 \inv[3370]/_0_  (.A(\inv_in[3370] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3371] ));
 sky130_fd_sc_hd__inv_2 \inv[3371]/_0_  (.A(\inv_in[3371] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3372] ));
 sky130_fd_sc_hd__inv_2 \inv[3372]/_0_  (.A(\inv_in[3372] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3373] ));
 sky130_fd_sc_hd__inv_2 \inv[3373]/_0_  (.A(\inv_in[3373] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3374] ));
 sky130_fd_sc_hd__inv_2 \inv[3374]/_0_  (.A(\inv_in[3374] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3375] ));
 sky130_fd_sc_hd__inv_2 \inv[3375]/_0_  (.A(\inv_in[3375] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3376] ));
 sky130_fd_sc_hd__inv_2 \inv[3376]/_0_  (.A(\inv_in[3376] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3377] ));
 sky130_fd_sc_hd__inv_2 \inv[3377]/_0_  (.A(\inv_in[3377] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3378] ));
 sky130_fd_sc_hd__inv_2 \inv[3378]/_0_  (.A(\inv_in[3378] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3379] ));
 sky130_fd_sc_hd__inv_2 \inv[3379]/_0_  (.A(\inv_in[3379] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3380] ));
 sky130_fd_sc_hd__inv_2 \inv[337]/_0_  (.A(\inv_in[337] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[338] ));
 sky130_fd_sc_hd__inv_2 \inv[3380]/_0_  (.A(\inv_in[3380] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3381] ));
 sky130_fd_sc_hd__inv_2 \inv[3381]/_0_  (.A(\inv_in[3381] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3382] ));
 sky130_fd_sc_hd__inv_2 \inv[3382]/_0_  (.A(\inv_in[3382] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3383] ));
 sky130_fd_sc_hd__inv_2 \inv[3383]/_0_  (.A(\inv_in[3383] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3384] ));
 sky130_fd_sc_hd__inv_2 \inv[3384]/_0_  (.A(\inv_in[3384] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3385] ));
 sky130_fd_sc_hd__inv_2 \inv[3385]/_0_  (.A(\inv_in[3385] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3386] ));
 sky130_fd_sc_hd__inv_2 \inv[3386]/_0_  (.A(\inv_in[3386] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3387] ));
 sky130_fd_sc_hd__inv_2 \inv[3387]/_0_  (.A(\inv_in[3387] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3388] ));
 sky130_fd_sc_hd__inv_2 \inv[3388]/_0_  (.A(\inv_in[3388] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3389] ));
 sky130_fd_sc_hd__inv_2 \inv[3389]/_0_  (.A(\inv_in[3389] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3390] ));
 sky130_fd_sc_hd__inv_2 \inv[338]/_0_  (.A(\inv_in[338] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[339] ));
 sky130_fd_sc_hd__inv_2 \inv[3390]/_0_  (.A(\inv_in[3390] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3391] ));
 sky130_fd_sc_hd__inv_2 \inv[3391]/_0_  (.A(\inv_in[3391] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3392] ));
 sky130_fd_sc_hd__inv_2 \inv[3392]/_0_  (.A(\inv_in[3392] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3393] ));
 sky130_fd_sc_hd__inv_2 \inv[3393]/_0_  (.A(\inv_in[3393] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3394] ));
 sky130_fd_sc_hd__inv_2 \inv[3394]/_0_  (.A(\inv_in[3394] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3395] ));
 sky130_fd_sc_hd__inv_2 \inv[3395]/_0_  (.A(\inv_in[3395] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3396] ));
 sky130_fd_sc_hd__inv_2 \inv[3396]/_0_  (.A(\inv_in[3396] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3397] ));
 sky130_fd_sc_hd__inv_2 \inv[3397]/_0_  (.A(\inv_in[3397] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3398] ));
 sky130_fd_sc_hd__inv_2 \inv[3398]/_0_  (.A(\inv_in[3398] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3399] ));
 sky130_fd_sc_hd__inv_2 \inv[3399]/_0_  (.A(\inv_in[3399] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3400] ));
 sky130_fd_sc_hd__inv_2 \inv[339]/_0_  (.A(\inv_in[339] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[340] ));
 sky130_fd_sc_hd__inv_2 \inv[33]/_0_  (.A(\inv_in[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[34] ));
 sky130_fd_sc_hd__inv_2 \inv[3400]/_0_  (.A(\inv_in[3400] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3401] ));
 sky130_fd_sc_hd__inv_2 \inv[3401]/_0_  (.A(\inv_in[3401] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3402] ));
 sky130_fd_sc_hd__inv_2 \inv[3402]/_0_  (.A(\inv_in[3402] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3403] ));
 sky130_fd_sc_hd__inv_2 \inv[3403]/_0_  (.A(\inv_in[3403] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3404] ));
 sky130_fd_sc_hd__inv_2 \inv[3404]/_0_  (.A(\inv_in[3404] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3405] ));
 sky130_fd_sc_hd__inv_2 \inv[3405]/_0_  (.A(\inv_in[3405] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3406] ));
 sky130_fd_sc_hd__inv_2 \inv[3406]/_0_  (.A(\inv_in[3406] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3407] ));
 sky130_fd_sc_hd__inv_2 \inv[3407]/_0_  (.A(\inv_in[3407] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3408] ));
 sky130_fd_sc_hd__inv_2 \inv[3408]/_0_  (.A(\inv_in[3408] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3409] ));
 sky130_fd_sc_hd__inv_2 \inv[3409]/_0_  (.A(\inv_in[3409] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3410] ));
 sky130_fd_sc_hd__inv_2 \inv[340]/_0_  (.A(\inv_in[340] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[341] ));
 sky130_fd_sc_hd__inv_2 \inv[3410]/_0_  (.A(\inv_in[3410] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3411] ));
 sky130_fd_sc_hd__inv_2 \inv[3411]/_0_  (.A(\inv_in[3411] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3412] ));
 sky130_fd_sc_hd__inv_2 \inv[3412]/_0_  (.A(\inv_in[3412] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3413] ));
 sky130_fd_sc_hd__inv_2 \inv[3413]/_0_  (.A(\inv_in[3413] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3414] ));
 sky130_fd_sc_hd__inv_2 \inv[3414]/_0_  (.A(\inv_in[3414] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3415] ));
 sky130_fd_sc_hd__inv_2 \inv[3415]/_0_  (.A(\inv_in[3415] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3416] ));
 sky130_fd_sc_hd__inv_2 \inv[3416]/_0_  (.A(\inv_in[3416] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3417] ));
 sky130_fd_sc_hd__inv_2 \inv[3417]/_0_  (.A(\inv_in[3417] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3418] ));
 sky130_fd_sc_hd__inv_2 \inv[3418]/_0_  (.A(\inv_in[3418] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3419] ));
 sky130_fd_sc_hd__inv_2 \inv[3419]/_0_  (.A(\inv_in[3419] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3420] ));
 sky130_fd_sc_hd__inv_2 \inv[341]/_0_  (.A(\inv_in[341] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[342] ));
 sky130_fd_sc_hd__inv_2 \inv[3420]/_0_  (.A(\inv_in[3420] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3421] ));
 sky130_fd_sc_hd__inv_2 \inv[3421]/_0_  (.A(\inv_in[3421] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3422] ));
 sky130_fd_sc_hd__inv_2 \inv[3422]/_0_  (.A(\inv_in[3422] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3423] ));
 sky130_fd_sc_hd__inv_2 \inv[3423]/_0_  (.A(\inv_in[3423] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3424] ));
 sky130_fd_sc_hd__inv_2 \inv[3424]/_0_  (.A(\inv_in[3424] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3425] ));
 sky130_fd_sc_hd__inv_2 \inv[3425]/_0_  (.A(\inv_in[3425] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3426] ));
 sky130_fd_sc_hd__inv_2 \inv[3426]/_0_  (.A(\inv_in[3426] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3427] ));
 sky130_fd_sc_hd__inv_2 \inv[3427]/_0_  (.A(\inv_in[3427] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3428] ));
 sky130_fd_sc_hd__inv_2 \inv[3428]/_0_  (.A(\inv_in[3428] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3429] ));
 sky130_fd_sc_hd__inv_2 \inv[3429]/_0_  (.A(\inv_in[3429] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3430] ));
 sky130_fd_sc_hd__inv_2 \inv[342]/_0_  (.A(\inv_in[342] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[343] ));
 sky130_fd_sc_hd__inv_2 \inv[3430]/_0_  (.A(\inv_in[3430] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3431] ));
 sky130_fd_sc_hd__inv_2 \inv[3431]/_0_  (.A(\inv_in[3431] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3432] ));
 sky130_fd_sc_hd__inv_2 \inv[3432]/_0_  (.A(\inv_in[3432] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3433] ));
 sky130_fd_sc_hd__inv_2 \inv[3433]/_0_  (.A(\inv_in[3433] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3434] ));
 sky130_fd_sc_hd__inv_2 \inv[3434]/_0_  (.A(\inv_in[3434] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3435] ));
 sky130_fd_sc_hd__inv_2 \inv[3435]/_0_  (.A(\inv_in[3435] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3436] ));
 sky130_fd_sc_hd__inv_2 \inv[3436]/_0_  (.A(\inv_in[3436] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3437] ));
 sky130_fd_sc_hd__inv_2 \inv[3437]/_0_  (.A(\inv_in[3437] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3438] ));
 sky130_fd_sc_hd__inv_2 \inv[3438]/_0_  (.A(\inv_in[3438] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3439] ));
 sky130_fd_sc_hd__inv_2 \inv[3439]/_0_  (.A(\inv_in[3439] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3440] ));
 sky130_fd_sc_hd__inv_2 \inv[343]/_0_  (.A(\inv_in[343] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[344] ));
 sky130_fd_sc_hd__inv_2 \inv[3440]/_0_  (.A(\inv_in[3440] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3441] ));
 sky130_fd_sc_hd__inv_2 \inv[3441]/_0_  (.A(\inv_in[3441] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3442] ));
 sky130_fd_sc_hd__inv_2 \inv[3442]/_0_  (.A(\inv_in[3442] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3443] ));
 sky130_fd_sc_hd__inv_2 \inv[3443]/_0_  (.A(\inv_in[3443] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3444] ));
 sky130_fd_sc_hd__inv_2 \inv[3444]/_0_  (.A(\inv_in[3444] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3445] ));
 sky130_fd_sc_hd__inv_2 \inv[3445]/_0_  (.A(\inv_in[3445] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3446] ));
 sky130_fd_sc_hd__inv_2 \inv[3446]/_0_  (.A(\inv_in[3446] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3447] ));
 sky130_fd_sc_hd__inv_2 \inv[3447]/_0_  (.A(\inv_in[3447] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3448] ));
 sky130_fd_sc_hd__inv_2 \inv[3448]/_0_  (.A(\inv_in[3448] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3449] ));
 sky130_fd_sc_hd__inv_2 \inv[3449]/_0_  (.A(\inv_in[3449] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3450] ));
 sky130_fd_sc_hd__inv_2 \inv[344]/_0_  (.A(\inv_in[344] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[345] ));
 sky130_fd_sc_hd__inv_2 \inv[3450]/_0_  (.A(\inv_in[3450] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3451] ));
 sky130_fd_sc_hd__inv_2 \inv[3451]/_0_  (.A(\inv_in[3451] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3452] ));
 sky130_fd_sc_hd__inv_2 \inv[3452]/_0_  (.A(\inv_in[3452] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3453] ));
 sky130_fd_sc_hd__inv_2 \inv[3453]/_0_  (.A(\inv_in[3453] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3454] ));
 sky130_fd_sc_hd__inv_2 \inv[3454]/_0_  (.A(\inv_in[3454] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3455] ));
 sky130_fd_sc_hd__inv_2 \inv[3455]/_0_  (.A(\inv_in[3455] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3456] ));
 sky130_fd_sc_hd__inv_2 \inv[3456]/_0_  (.A(\inv_in[3456] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3457] ));
 sky130_fd_sc_hd__inv_2 \inv[3457]/_0_  (.A(\inv_in[3457] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3458] ));
 sky130_fd_sc_hd__inv_2 \inv[3458]/_0_  (.A(\inv_in[3458] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3459] ));
 sky130_fd_sc_hd__inv_2 \inv[3459]/_0_  (.A(\inv_in[3459] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3460] ));
 sky130_fd_sc_hd__inv_2 \inv[345]/_0_  (.A(\inv_in[345] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[346] ));
 sky130_fd_sc_hd__inv_2 \inv[3460]/_0_  (.A(\inv_in[3460] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3461] ));
 sky130_fd_sc_hd__inv_2 \inv[3461]/_0_  (.A(\inv_in[3461] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3462] ));
 sky130_fd_sc_hd__inv_2 \inv[3462]/_0_  (.A(\inv_in[3462] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3463] ));
 sky130_fd_sc_hd__inv_2 \inv[3463]/_0_  (.A(\inv_in[3463] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3464] ));
 sky130_fd_sc_hd__inv_2 \inv[3464]/_0_  (.A(\inv_in[3464] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3465] ));
 sky130_fd_sc_hd__inv_2 \inv[3465]/_0_  (.A(\inv_in[3465] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3466] ));
 sky130_fd_sc_hd__inv_2 \inv[3466]/_0_  (.A(\inv_in[3466] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3467] ));
 sky130_fd_sc_hd__inv_2 \inv[3467]/_0_  (.A(\inv_in[3467] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3468] ));
 sky130_fd_sc_hd__inv_2 \inv[3468]/_0_  (.A(\inv_in[3468] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3469] ));
 sky130_fd_sc_hd__inv_2 \inv[3469]/_0_  (.A(\inv_in[3469] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3470] ));
 sky130_fd_sc_hd__inv_2 \inv[346]/_0_  (.A(\inv_in[346] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[347] ));
 sky130_fd_sc_hd__inv_2 \inv[3470]/_0_  (.A(\inv_in[3470] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3471] ));
 sky130_fd_sc_hd__inv_2 \inv[3471]/_0_  (.A(\inv_in[3471] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3472] ));
 sky130_fd_sc_hd__inv_2 \inv[3472]/_0_  (.A(\inv_in[3472] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3473] ));
 sky130_fd_sc_hd__inv_2 \inv[3473]/_0_  (.A(\inv_in[3473] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3474] ));
 sky130_fd_sc_hd__inv_2 \inv[3474]/_0_  (.A(\inv_in[3474] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3475] ));
 sky130_fd_sc_hd__inv_2 \inv[3475]/_0_  (.A(\inv_in[3475] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3476] ));
 sky130_fd_sc_hd__inv_2 \inv[3476]/_0_  (.A(\inv_in[3476] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3477] ));
 sky130_fd_sc_hd__inv_2 \inv[3477]/_0_  (.A(\inv_in[3477] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3478] ));
 sky130_fd_sc_hd__inv_2 \inv[3478]/_0_  (.A(\inv_in[3478] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3479] ));
 sky130_fd_sc_hd__inv_2 \inv[3479]/_0_  (.A(\inv_in[3479] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3480] ));
 sky130_fd_sc_hd__inv_2 \inv[347]/_0_  (.A(\inv_in[347] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[348] ));
 sky130_fd_sc_hd__inv_2 \inv[3480]/_0_  (.A(\inv_in[3480] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3481] ));
 sky130_fd_sc_hd__inv_2 \inv[3481]/_0_  (.A(\inv_in[3481] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3482] ));
 sky130_fd_sc_hd__inv_2 \inv[3482]/_0_  (.A(\inv_in[3482] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3483] ));
 sky130_fd_sc_hd__inv_2 \inv[3483]/_0_  (.A(\inv_in[3483] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3484] ));
 sky130_fd_sc_hd__inv_2 \inv[3484]/_0_  (.A(\inv_in[3484] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3485] ));
 sky130_fd_sc_hd__inv_2 \inv[3485]/_0_  (.A(\inv_in[3485] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3486] ));
 sky130_fd_sc_hd__inv_2 \inv[3486]/_0_  (.A(\inv_in[3486] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3487] ));
 sky130_fd_sc_hd__inv_2 \inv[3487]/_0_  (.A(\inv_in[3487] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3488] ));
 sky130_fd_sc_hd__inv_2 \inv[3488]/_0_  (.A(\inv_in[3488] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3489] ));
 sky130_fd_sc_hd__inv_2 \inv[3489]/_0_  (.A(\inv_in[3489] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3490] ));
 sky130_fd_sc_hd__inv_2 \inv[348]/_0_  (.A(\inv_in[348] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[349] ));
 sky130_fd_sc_hd__inv_2 \inv[3490]/_0_  (.A(\inv_in[3490] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3491] ));
 sky130_fd_sc_hd__inv_2 \inv[3491]/_0_  (.A(\inv_in[3491] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3492] ));
 sky130_fd_sc_hd__inv_2 \inv[3492]/_0_  (.A(\inv_in[3492] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3493] ));
 sky130_fd_sc_hd__inv_2 \inv[3493]/_0_  (.A(\inv_in[3493] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3494] ));
 sky130_fd_sc_hd__inv_2 \inv[3494]/_0_  (.A(\inv_in[3494] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3495] ));
 sky130_fd_sc_hd__inv_2 \inv[3495]/_0_  (.A(\inv_in[3495] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3496] ));
 sky130_fd_sc_hd__inv_2 \inv[3496]/_0_  (.A(\inv_in[3496] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3497] ));
 sky130_fd_sc_hd__inv_2 \inv[3497]/_0_  (.A(\inv_in[3497] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3498] ));
 sky130_fd_sc_hd__inv_2 \inv[3498]/_0_  (.A(\inv_in[3498] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3499] ));
 sky130_fd_sc_hd__inv_2 \inv[3499]/_0_  (.A(\inv_in[3499] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3500] ));
 sky130_fd_sc_hd__inv_2 \inv[349]/_0_  (.A(\inv_in[349] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[350] ));
 sky130_fd_sc_hd__inv_2 \inv[34]/_0_  (.A(\inv_in[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[35] ));
 sky130_fd_sc_hd__inv_2 \inv[3500]/_0_  (.A(\inv_in[3500] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3501] ));
 sky130_fd_sc_hd__inv_2 \inv[3501]/_0_  (.A(\inv_in[3501] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3502] ));
 sky130_fd_sc_hd__inv_2 \inv[3502]/_0_  (.A(\inv_in[3502] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3503] ));
 sky130_fd_sc_hd__inv_2 \inv[3503]/_0_  (.A(\inv_in[3503] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3504] ));
 sky130_fd_sc_hd__inv_2 \inv[3504]/_0_  (.A(\inv_in[3504] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3505] ));
 sky130_fd_sc_hd__inv_2 \inv[3505]/_0_  (.A(\inv_in[3505] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3506] ));
 sky130_fd_sc_hd__inv_2 \inv[3506]/_0_  (.A(\inv_in[3506] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3507] ));
 sky130_fd_sc_hd__inv_2 \inv[3507]/_0_  (.A(\inv_in[3507] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3508] ));
 sky130_fd_sc_hd__inv_2 \inv[3508]/_0_  (.A(\inv_in[3508] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3509] ));
 sky130_fd_sc_hd__inv_2 \inv[3509]/_0_  (.A(\inv_in[3509] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3510] ));
 sky130_fd_sc_hd__inv_2 \inv[350]/_0_  (.A(\inv_in[350] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[351] ));
 sky130_fd_sc_hd__inv_2 \inv[3510]/_0_  (.A(\inv_in[3510] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3511] ));
 sky130_fd_sc_hd__inv_2 \inv[3511]/_0_  (.A(\inv_in[3511] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3512] ));
 sky130_fd_sc_hd__inv_2 \inv[3512]/_0_  (.A(\inv_in[3512] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3513] ));
 sky130_fd_sc_hd__inv_2 \inv[3513]/_0_  (.A(\inv_in[3513] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3514] ));
 sky130_fd_sc_hd__inv_2 \inv[3514]/_0_  (.A(\inv_in[3514] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3515] ));
 sky130_fd_sc_hd__inv_2 \inv[3515]/_0_  (.A(\inv_in[3515] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3516] ));
 sky130_fd_sc_hd__inv_2 \inv[3516]/_0_  (.A(\inv_in[3516] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3517] ));
 sky130_fd_sc_hd__inv_2 \inv[3517]/_0_  (.A(\inv_in[3517] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3518] ));
 sky130_fd_sc_hd__inv_2 \inv[3518]/_0_  (.A(\inv_in[3518] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3519] ));
 sky130_fd_sc_hd__inv_2 \inv[3519]/_0_  (.A(\inv_in[3519] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3520] ));
 sky130_fd_sc_hd__inv_2 \inv[351]/_0_  (.A(\inv_in[351] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[352] ));
 sky130_fd_sc_hd__inv_2 \inv[3520]/_0_  (.A(\inv_in[3520] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3521] ));
 sky130_fd_sc_hd__inv_2 \inv[3521]/_0_  (.A(\inv_in[3521] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3522] ));
 sky130_fd_sc_hd__inv_2 \inv[3522]/_0_  (.A(\inv_in[3522] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3523] ));
 sky130_fd_sc_hd__inv_2 \inv[3523]/_0_  (.A(\inv_in[3523] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3524] ));
 sky130_fd_sc_hd__inv_2 \inv[3524]/_0_  (.A(\inv_in[3524] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3525] ));
 sky130_fd_sc_hd__inv_2 \inv[3525]/_0_  (.A(\inv_in[3525] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3526] ));
 sky130_fd_sc_hd__inv_2 \inv[3526]/_0_  (.A(\inv_in[3526] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3527] ));
 sky130_fd_sc_hd__inv_2 \inv[3527]/_0_  (.A(\inv_in[3527] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3528] ));
 sky130_fd_sc_hd__inv_2 \inv[3528]/_0_  (.A(\inv_in[3528] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3529] ));
 sky130_fd_sc_hd__inv_2 \inv[3529]/_0_  (.A(\inv_in[3529] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3530] ));
 sky130_fd_sc_hd__inv_2 \inv[352]/_0_  (.A(\inv_in[352] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[353] ));
 sky130_fd_sc_hd__inv_2 \inv[3530]/_0_  (.A(\inv_in[3530] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3531] ));
 sky130_fd_sc_hd__inv_2 \inv[3531]/_0_  (.A(\inv_in[3531] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3532] ));
 sky130_fd_sc_hd__inv_2 \inv[3532]/_0_  (.A(\inv_in[3532] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3533] ));
 sky130_fd_sc_hd__inv_2 \inv[3533]/_0_  (.A(\inv_in[3533] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3534] ));
 sky130_fd_sc_hd__inv_2 \inv[3534]/_0_  (.A(\inv_in[3534] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3535] ));
 sky130_fd_sc_hd__inv_2 \inv[3535]/_0_  (.A(\inv_in[3535] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3536] ));
 sky130_fd_sc_hd__inv_2 \inv[3536]/_0_  (.A(\inv_in[3536] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3537] ));
 sky130_fd_sc_hd__inv_2 \inv[3537]/_0_  (.A(\inv_in[3537] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3538] ));
 sky130_fd_sc_hd__inv_2 \inv[3538]/_0_  (.A(\inv_in[3538] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3539] ));
 sky130_fd_sc_hd__inv_2 \inv[3539]/_0_  (.A(\inv_in[3539] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3540] ));
 sky130_fd_sc_hd__inv_2 \inv[353]/_0_  (.A(\inv_in[353] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[354] ));
 sky130_fd_sc_hd__inv_2 \inv[3540]/_0_  (.A(\inv_in[3540] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3541] ));
 sky130_fd_sc_hd__inv_2 \inv[3541]/_0_  (.A(\inv_in[3541] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3542] ));
 sky130_fd_sc_hd__inv_2 \inv[3542]/_0_  (.A(\inv_in[3542] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3543] ));
 sky130_fd_sc_hd__inv_2 \inv[3543]/_0_  (.A(\inv_in[3543] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3544] ));
 sky130_fd_sc_hd__inv_2 \inv[3544]/_0_  (.A(\inv_in[3544] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3545] ));
 sky130_fd_sc_hd__inv_2 \inv[3545]/_0_  (.A(\inv_in[3545] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3546] ));
 sky130_fd_sc_hd__inv_2 \inv[3546]/_0_  (.A(\inv_in[3546] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3547] ));
 sky130_fd_sc_hd__inv_2 \inv[3547]/_0_  (.A(\inv_in[3547] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3548] ));
 sky130_fd_sc_hd__inv_2 \inv[3548]/_0_  (.A(\inv_in[3548] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3549] ));
 sky130_fd_sc_hd__inv_2 \inv[3549]/_0_  (.A(\inv_in[3549] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3550] ));
 sky130_fd_sc_hd__inv_2 \inv[354]/_0_  (.A(\inv_in[354] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[355] ));
 sky130_fd_sc_hd__inv_2 \inv[3550]/_0_  (.A(\inv_in[3550] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3551] ));
 sky130_fd_sc_hd__inv_2 \inv[3551]/_0_  (.A(\inv_in[3551] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3552] ));
 sky130_fd_sc_hd__inv_2 \inv[3552]/_0_  (.A(\inv_in[3552] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3553] ));
 sky130_fd_sc_hd__inv_2 \inv[3553]/_0_  (.A(\inv_in[3553] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3554] ));
 sky130_fd_sc_hd__inv_2 \inv[3554]/_0_  (.A(\inv_in[3554] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3555] ));
 sky130_fd_sc_hd__inv_2 \inv[3555]/_0_  (.A(\inv_in[3555] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3556] ));
 sky130_fd_sc_hd__inv_2 \inv[3556]/_0_  (.A(\inv_in[3556] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3557] ));
 sky130_fd_sc_hd__inv_2 \inv[3557]/_0_  (.A(\inv_in[3557] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3558] ));
 sky130_fd_sc_hd__inv_2 \inv[3558]/_0_  (.A(\inv_in[3558] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3559] ));
 sky130_fd_sc_hd__inv_2 \inv[3559]/_0_  (.A(\inv_in[3559] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3560] ));
 sky130_fd_sc_hd__inv_2 \inv[355]/_0_  (.A(\inv_in[355] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[356] ));
 sky130_fd_sc_hd__inv_2 \inv[3560]/_0_  (.A(\inv_in[3560] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3561] ));
 sky130_fd_sc_hd__inv_2 \inv[3561]/_0_  (.A(\inv_in[3561] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3562] ));
 sky130_fd_sc_hd__inv_2 \inv[3562]/_0_  (.A(\inv_in[3562] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3563] ));
 sky130_fd_sc_hd__inv_2 \inv[3563]/_0_  (.A(\inv_in[3563] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3564] ));
 sky130_fd_sc_hd__inv_2 \inv[3564]/_0_  (.A(\inv_in[3564] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3565] ));
 sky130_fd_sc_hd__inv_2 \inv[3565]/_0_  (.A(\inv_in[3565] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3566] ));
 sky130_fd_sc_hd__inv_2 \inv[3566]/_0_  (.A(\inv_in[3566] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3567] ));
 sky130_fd_sc_hd__inv_2 \inv[3567]/_0_  (.A(\inv_in[3567] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3568] ));
 sky130_fd_sc_hd__inv_2 \inv[3568]/_0_  (.A(\inv_in[3568] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3569] ));
 sky130_fd_sc_hd__inv_2 \inv[3569]/_0_  (.A(\inv_in[3569] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3570] ));
 sky130_fd_sc_hd__inv_2 \inv[356]/_0_  (.A(\inv_in[356] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[357] ));
 sky130_fd_sc_hd__inv_2 \inv[3570]/_0_  (.A(\inv_in[3570] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3571] ));
 sky130_fd_sc_hd__inv_2 \inv[3571]/_0_  (.A(\inv_in[3571] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3572] ));
 sky130_fd_sc_hd__inv_2 \inv[3572]/_0_  (.A(\inv_in[3572] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3573] ));
 sky130_fd_sc_hd__inv_2 \inv[3573]/_0_  (.A(\inv_in[3573] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3574] ));
 sky130_fd_sc_hd__inv_2 \inv[3574]/_0_  (.A(\inv_in[3574] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3575] ));
 sky130_fd_sc_hd__inv_2 \inv[3575]/_0_  (.A(\inv_in[3575] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3576] ));
 sky130_fd_sc_hd__inv_2 \inv[3576]/_0_  (.A(\inv_in[3576] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3577] ));
 sky130_fd_sc_hd__inv_2 \inv[3577]/_0_  (.A(\inv_in[3577] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3578] ));
 sky130_fd_sc_hd__inv_2 \inv[3578]/_0_  (.A(\inv_in[3578] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3579] ));
 sky130_fd_sc_hd__inv_2 \inv[3579]/_0_  (.A(\inv_in[3579] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3580] ));
 sky130_fd_sc_hd__inv_2 \inv[357]/_0_  (.A(\inv_in[357] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[358] ));
 sky130_fd_sc_hd__inv_2 \inv[3580]/_0_  (.A(\inv_in[3580] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3581] ));
 sky130_fd_sc_hd__inv_2 \inv[3581]/_0_  (.A(\inv_in[3581] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3582] ));
 sky130_fd_sc_hd__inv_2 \inv[3582]/_0_  (.A(\inv_in[3582] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3583] ));
 sky130_fd_sc_hd__inv_2 \inv[3583]/_0_  (.A(\inv_in[3583] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3584] ));
 sky130_fd_sc_hd__inv_2 \inv[3584]/_0_  (.A(\inv_in[3584] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3585] ));
 sky130_fd_sc_hd__inv_2 \inv[3585]/_0_  (.A(\inv_in[3585] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3586] ));
 sky130_fd_sc_hd__inv_2 \inv[3586]/_0_  (.A(\inv_in[3586] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3587] ));
 sky130_fd_sc_hd__inv_2 \inv[3587]/_0_  (.A(\inv_in[3587] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3588] ));
 sky130_fd_sc_hd__inv_2 \inv[3588]/_0_  (.A(\inv_in[3588] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3589] ));
 sky130_fd_sc_hd__inv_2 \inv[3589]/_0_  (.A(\inv_in[3589] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3590] ));
 sky130_fd_sc_hd__inv_2 \inv[358]/_0_  (.A(\inv_in[358] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[359] ));
 sky130_fd_sc_hd__inv_2 \inv[3590]/_0_  (.A(\inv_in[3590] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3591] ));
 sky130_fd_sc_hd__inv_2 \inv[3591]/_0_  (.A(\inv_in[3591] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3592] ));
 sky130_fd_sc_hd__inv_2 \inv[3592]/_0_  (.A(\inv_in[3592] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3593] ));
 sky130_fd_sc_hd__inv_2 \inv[3593]/_0_  (.A(\inv_in[3593] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3594] ));
 sky130_fd_sc_hd__inv_2 \inv[3594]/_0_  (.A(\inv_in[3594] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3595] ));
 sky130_fd_sc_hd__inv_2 \inv[3595]/_0_  (.A(\inv_in[3595] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3596] ));
 sky130_fd_sc_hd__inv_2 \inv[3596]/_0_  (.A(\inv_in[3596] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3597] ));
 sky130_fd_sc_hd__inv_2 \inv[3597]/_0_  (.A(\inv_in[3597] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3598] ));
 sky130_fd_sc_hd__inv_2 \inv[3598]/_0_  (.A(\inv_in[3598] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3599] ));
 sky130_fd_sc_hd__inv_2 \inv[3599]/_0_  (.A(\inv_in[3599] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3600] ));
 sky130_fd_sc_hd__inv_2 \inv[359]/_0_  (.A(\inv_in[359] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[360] ));
 sky130_fd_sc_hd__inv_2 \inv[35]/_0_  (.A(\inv_in[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[36] ));
 sky130_fd_sc_hd__inv_2 \inv[3600]/_0_  (.A(\inv_in[3600] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3601] ));
 sky130_fd_sc_hd__inv_2 \inv[3601]/_0_  (.A(\inv_in[3601] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3602] ));
 sky130_fd_sc_hd__inv_2 \inv[3602]/_0_  (.A(\inv_in[3602] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3603] ));
 sky130_fd_sc_hd__inv_2 \inv[3603]/_0_  (.A(\inv_in[3603] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3604] ));
 sky130_fd_sc_hd__inv_2 \inv[3604]/_0_  (.A(\inv_in[3604] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3605] ));
 sky130_fd_sc_hd__inv_2 \inv[3605]/_0_  (.A(\inv_in[3605] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3606] ));
 sky130_fd_sc_hd__inv_2 \inv[3606]/_0_  (.A(\inv_in[3606] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3607] ));
 sky130_fd_sc_hd__inv_2 \inv[3607]/_0_  (.A(\inv_in[3607] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3608] ));
 sky130_fd_sc_hd__inv_2 \inv[3608]/_0_  (.A(\inv_in[3608] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3609] ));
 sky130_fd_sc_hd__inv_2 \inv[3609]/_0_  (.A(\inv_in[3609] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3610] ));
 sky130_fd_sc_hd__inv_2 \inv[360]/_0_  (.A(\inv_in[360] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[361] ));
 sky130_fd_sc_hd__inv_2 \inv[3610]/_0_  (.A(\inv_in[3610] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3611] ));
 sky130_fd_sc_hd__inv_2 \inv[3611]/_0_  (.A(\inv_in[3611] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3612] ));
 sky130_fd_sc_hd__inv_2 \inv[3612]/_0_  (.A(\inv_in[3612] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3613] ));
 sky130_fd_sc_hd__inv_2 \inv[3613]/_0_  (.A(\inv_in[3613] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3614] ));
 sky130_fd_sc_hd__inv_2 \inv[3614]/_0_  (.A(\inv_in[3614] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3615] ));
 sky130_fd_sc_hd__inv_2 \inv[3615]/_0_  (.A(\inv_in[3615] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3616] ));
 sky130_fd_sc_hd__inv_2 \inv[3616]/_0_  (.A(\inv_in[3616] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3617] ));
 sky130_fd_sc_hd__inv_2 \inv[3617]/_0_  (.A(\inv_in[3617] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3618] ));
 sky130_fd_sc_hd__inv_2 \inv[3618]/_0_  (.A(\inv_in[3618] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3619] ));
 sky130_fd_sc_hd__inv_2 \inv[3619]/_0_  (.A(\inv_in[3619] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3620] ));
 sky130_fd_sc_hd__inv_2 \inv[361]/_0_  (.A(\inv_in[361] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[362] ));
 sky130_fd_sc_hd__inv_2 \inv[3620]/_0_  (.A(\inv_in[3620] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3621] ));
 sky130_fd_sc_hd__inv_2 \inv[3621]/_0_  (.A(\inv_in[3621] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3622] ));
 sky130_fd_sc_hd__inv_2 \inv[3622]/_0_  (.A(\inv_in[3622] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3623] ));
 sky130_fd_sc_hd__inv_2 \inv[3623]/_0_  (.A(\inv_in[3623] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3624] ));
 sky130_fd_sc_hd__inv_2 \inv[3624]/_0_  (.A(\inv_in[3624] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3625] ));
 sky130_fd_sc_hd__inv_2 \inv[3625]/_0_  (.A(\inv_in[3625] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3626] ));
 sky130_fd_sc_hd__inv_2 \inv[3626]/_0_  (.A(\inv_in[3626] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3627] ));
 sky130_fd_sc_hd__inv_2 \inv[3627]/_0_  (.A(\inv_in[3627] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3628] ));
 sky130_fd_sc_hd__inv_2 \inv[3628]/_0_  (.A(\inv_in[3628] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3629] ));
 sky130_fd_sc_hd__inv_2 \inv[3629]/_0_  (.A(\inv_in[3629] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3630] ));
 sky130_fd_sc_hd__inv_2 \inv[362]/_0_  (.A(\inv_in[362] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[363] ));
 sky130_fd_sc_hd__inv_2 \inv[3630]/_0_  (.A(\inv_in[3630] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3631] ));
 sky130_fd_sc_hd__inv_2 \inv[3631]/_0_  (.A(\inv_in[3631] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3632] ));
 sky130_fd_sc_hd__inv_2 \inv[3632]/_0_  (.A(\inv_in[3632] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3633] ));
 sky130_fd_sc_hd__inv_2 \inv[3633]/_0_  (.A(\inv_in[3633] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3634] ));
 sky130_fd_sc_hd__inv_2 \inv[3634]/_0_  (.A(\inv_in[3634] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3635] ));
 sky130_fd_sc_hd__inv_2 \inv[3635]/_0_  (.A(\inv_in[3635] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3636] ));
 sky130_fd_sc_hd__inv_2 \inv[3636]/_0_  (.A(\inv_in[3636] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3637] ));
 sky130_fd_sc_hd__inv_2 \inv[3637]/_0_  (.A(\inv_in[3637] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3638] ));
 sky130_fd_sc_hd__inv_2 \inv[3638]/_0_  (.A(\inv_in[3638] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3639] ));
 sky130_fd_sc_hd__inv_2 \inv[3639]/_0_  (.A(\inv_in[3639] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3640] ));
 sky130_fd_sc_hd__inv_2 \inv[363]/_0_  (.A(\inv_in[363] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[364] ));
 sky130_fd_sc_hd__inv_2 \inv[3640]/_0_  (.A(\inv_in[3640] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3641] ));
 sky130_fd_sc_hd__inv_2 \inv[3641]/_0_  (.A(\inv_in[3641] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3642] ));
 sky130_fd_sc_hd__inv_2 \inv[3642]/_0_  (.A(\inv_in[3642] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3643] ));
 sky130_fd_sc_hd__inv_2 \inv[3643]/_0_  (.A(\inv_in[3643] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3644] ));
 sky130_fd_sc_hd__inv_2 \inv[3644]/_0_  (.A(\inv_in[3644] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3645] ));
 sky130_fd_sc_hd__inv_2 \inv[3645]/_0_  (.A(\inv_in[3645] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3646] ));
 sky130_fd_sc_hd__inv_2 \inv[3646]/_0_  (.A(\inv_in[3646] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3647] ));
 sky130_fd_sc_hd__inv_2 \inv[3647]/_0_  (.A(\inv_in[3647] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3648] ));
 sky130_fd_sc_hd__inv_2 \inv[3648]/_0_  (.A(\inv_in[3648] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3649] ));
 sky130_fd_sc_hd__inv_2 \inv[3649]/_0_  (.A(\inv_in[3649] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3650] ));
 sky130_fd_sc_hd__inv_2 \inv[364]/_0_  (.A(\inv_in[364] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[365] ));
 sky130_fd_sc_hd__inv_2 \inv[3650]/_0_  (.A(\inv_in[3650] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3651] ));
 sky130_fd_sc_hd__inv_2 \inv[3651]/_0_  (.A(\inv_in[3651] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3652] ));
 sky130_fd_sc_hd__inv_2 \inv[3652]/_0_  (.A(\inv_in[3652] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3653] ));
 sky130_fd_sc_hd__inv_2 \inv[3653]/_0_  (.A(\inv_in[3653] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3654] ));
 sky130_fd_sc_hd__inv_2 \inv[3654]/_0_  (.A(\inv_in[3654] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3655] ));
 sky130_fd_sc_hd__inv_2 \inv[3655]/_0_  (.A(\inv_in[3655] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3656] ));
 sky130_fd_sc_hd__inv_2 \inv[3656]/_0_  (.A(\inv_in[3656] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3657] ));
 sky130_fd_sc_hd__inv_2 \inv[3657]/_0_  (.A(\inv_in[3657] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3658] ));
 sky130_fd_sc_hd__inv_2 \inv[3658]/_0_  (.A(\inv_in[3658] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3659] ));
 sky130_fd_sc_hd__inv_2 \inv[3659]/_0_  (.A(\inv_in[3659] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3660] ));
 sky130_fd_sc_hd__inv_2 \inv[365]/_0_  (.A(\inv_in[365] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[366] ));
 sky130_fd_sc_hd__inv_2 \inv[3660]/_0_  (.A(\inv_in[3660] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3661] ));
 sky130_fd_sc_hd__inv_2 \inv[3661]/_0_  (.A(\inv_in[3661] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3662] ));
 sky130_fd_sc_hd__inv_2 \inv[3662]/_0_  (.A(\inv_in[3662] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3663] ));
 sky130_fd_sc_hd__inv_2 \inv[3663]/_0_  (.A(\inv_in[3663] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3664] ));
 sky130_fd_sc_hd__inv_2 \inv[3664]/_0_  (.A(\inv_in[3664] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3665] ));
 sky130_fd_sc_hd__inv_2 \inv[3665]/_0_  (.A(\inv_in[3665] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3666] ));
 sky130_fd_sc_hd__inv_2 \inv[3666]/_0_  (.A(\inv_in[3666] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3667] ));
 sky130_fd_sc_hd__inv_2 \inv[3667]/_0_  (.A(\inv_in[3667] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3668] ));
 sky130_fd_sc_hd__inv_2 \inv[3668]/_0_  (.A(\inv_in[3668] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3669] ));
 sky130_fd_sc_hd__inv_2 \inv[3669]/_0_  (.A(\inv_in[3669] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3670] ));
 sky130_fd_sc_hd__inv_2 \inv[366]/_0_  (.A(\inv_in[366] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[367] ));
 sky130_fd_sc_hd__inv_2 \inv[3670]/_0_  (.A(\inv_in[3670] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3671] ));
 sky130_fd_sc_hd__inv_2 \inv[3671]/_0_  (.A(\inv_in[3671] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3672] ));
 sky130_fd_sc_hd__inv_2 \inv[3672]/_0_  (.A(\inv_in[3672] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3673] ));
 sky130_fd_sc_hd__inv_2 \inv[3673]/_0_  (.A(\inv_in[3673] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3674] ));
 sky130_fd_sc_hd__inv_2 \inv[3674]/_0_  (.A(\inv_in[3674] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3675] ));
 sky130_fd_sc_hd__inv_2 \inv[3675]/_0_  (.A(\inv_in[3675] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3676] ));
 sky130_fd_sc_hd__inv_2 \inv[3676]/_0_  (.A(\inv_in[3676] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3677] ));
 sky130_fd_sc_hd__inv_2 \inv[3677]/_0_  (.A(\inv_in[3677] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3678] ));
 sky130_fd_sc_hd__inv_2 \inv[3678]/_0_  (.A(\inv_in[3678] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3679] ));
 sky130_fd_sc_hd__inv_2 \inv[3679]/_0_  (.A(\inv_in[3679] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3680] ));
 sky130_fd_sc_hd__inv_2 \inv[367]/_0_  (.A(\inv_in[367] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[368] ));
 sky130_fd_sc_hd__inv_2 \inv[3680]/_0_  (.A(\inv_in[3680] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3681] ));
 sky130_fd_sc_hd__inv_2 \inv[3681]/_0_  (.A(\inv_in[3681] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3682] ));
 sky130_fd_sc_hd__inv_2 \inv[3682]/_0_  (.A(\inv_in[3682] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3683] ));
 sky130_fd_sc_hd__inv_2 \inv[3683]/_0_  (.A(\inv_in[3683] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3684] ));
 sky130_fd_sc_hd__inv_2 \inv[3684]/_0_  (.A(\inv_in[3684] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3685] ));
 sky130_fd_sc_hd__inv_2 \inv[3685]/_0_  (.A(\inv_in[3685] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3686] ));
 sky130_fd_sc_hd__inv_2 \inv[3686]/_0_  (.A(\inv_in[3686] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3687] ));
 sky130_fd_sc_hd__inv_2 \inv[3687]/_0_  (.A(\inv_in[3687] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3688] ));
 sky130_fd_sc_hd__inv_2 \inv[3688]/_0_  (.A(\inv_in[3688] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3689] ));
 sky130_fd_sc_hd__inv_2 \inv[3689]/_0_  (.A(\inv_in[3689] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3690] ));
 sky130_fd_sc_hd__inv_2 \inv[368]/_0_  (.A(\inv_in[368] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[369] ));
 sky130_fd_sc_hd__inv_2 \inv[3690]/_0_  (.A(\inv_in[3690] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3691] ));
 sky130_fd_sc_hd__inv_2 \inv[3691]/_0_  (.A(\inv_in[3691] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3692] ));
 sky130_fd_sc_hd__inv_2 \inv[3692]/_0_  (.A(\inv_in[3692] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3693] ));
 sky130_fd_sc_hd__inv_2 \inv[3693]/_0_  (.A(\inv_in[3693] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3694] ));
 sky130_fd_sc_hd__inv_2 \inv[3694]/_0_  (.A(\inv_in[3694] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3695] ));
 sky130_fd_sc_hd__inv_2 \inv[3695]/_0_  (.A(\inv_in[3695] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3696] ));
 sky130_fd_sc_hd__inv_2 \inv[3696]/_0_  (.A(\inv_in[3696] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3697] ));
 sky130_fd_sc_hd__inv_2 \inv[3697]/_0_  (.A(\inv_in[3697] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3698] ));
 sky130_fd_sc_hd__inv_2 \inv[3698]/_0_  (.A(\inv_in[3698] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3699] ));
 sky130_fd_sc_hd__inv_2 \inv[3699]/_0_  (.A(\inv_in[3699] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3700] ));
 sky130_fd_sc_hd__inv_2 \inv[369]/_0_  (.A(\inv_in[369] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[370] ));
 sky130_fd_sc_hd__inv_2 \inv[36]/_0_  (.A(\inv_in[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[37] ));
 sky130_fd_sc_hd__inv_2 \inv[3700]/_0_  (.A(\inv_in[3700] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3701] ));
 sky130_fd_sc_hd__inv_2 \inv[3701]/_0_  (.A(\inv_in[3701] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3702] ));
 sky130_fd_sc_hd__inv_2 \inv[3702]/_0_  (.A(\inv_in[3702] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3703] ));
 sky130_fd_sc_hd__inv_2 \inv[3703]/_0_  (.A(\inv_in[3703] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3704] ));
 sky130_fd_sc_hd__inv_2 \inv[3704]/_0_  (.A(\inv_in[3704] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3705] ));
 sky130_fd_sc_hd__inv_2 \inv[3705]/_0_  (.A(\inv_in[3705] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3706] ));
 sky130_fd_sc_hd__inv_2 \inv[3706]/_0_  (.A(\inv_in[3706] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3707] ));
 sky130_fd_sc_hd__inv_2 \inv[3707]/_0_  (.A(\inv_in[3707] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3708] ));
 sky130_fd_sc_hd__inv_2 \inv[3708]/_0_  (.A(\inv_in[3708] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3709] ));
 sky130_fd_sc_hd__inv_2 \inv[3709]/_0_  (.A(\inv_in[3709] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3710] ));
 sky130_fd_sc_hd__inv_2 \inv[370]/_0_  (.A(\inv_in[370] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[371] ));
 sky130_fd_sc_hd__inv_2 \inv[3710]/_0_  (.A(\inv_in[3710] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3711] ));
 sky130_fd_sc_hd__inv_2 \inv[3711]/_0_  (.A(\inv_in[3711] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3712] ));
 sky130_fd_sc_hd__inv_2 \inv[3712]/_0_  (.A(\inv_in[3712] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3713] ));
 sky130_fd_sc_hd__inv_2 \inv[3713]/_0_  (.A(\inv_in[3713] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3714] ));
 sky130_fd_sc_hd__inv_2 \inv[3714]/_0_  (.A(\inv_in[3714] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3715] ));
 sky130_fd_sc_hd__inv_2 \inv[3715]/_0_  (.A(\inv_in[3715] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3716] ));
 sky130_fd_sc_hd__inv_2 \inv[3716]/_0_  (.A(\inv_in[3716] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3717] ));
 sky130_fd_sc_hd__inv_2 \inv[3717]/_0_  (.A(\inv_in[3717] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3718] ));
 sky130_fd_sc_hd__inv_2 \inv[3718]/_0_  (.A(\inv_in[3718] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3719] ));
 sky130_fd_sc_hd__inv_2 \inv[3719]/_0_  (.A(\inv_in[3719] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3720] ));
 sky130_fd_sc_hd__inv_2 \inv[371]/_0_  (.A(\inv_in[371] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[372] ));
 sky130_fd_sc_hd__inv_2 \inv[3720]/_0_  (.A(\inv_in[3720] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3721] ));
 sky130_fd_sc_hd__inv_2 \inv[3721]/_0_  (.A(\inv_in[3721] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3722] ));
 sky130_fd_sc_hd__inv_2 \inv[3722]/_0_  (.A(\inv_in[3722] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3723] ));
 sky130_fd_sc_hd__inv_2 \inv[3723]/_0_  (.A(\inv_in[3723] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3724] ));
 sky130_fd_sc_hd__inv_2 \inv[3724]/_0_  (.A(\inv_in[3724] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3725] ));
 sky130_fd_sc_hd__inv_2 \inv[3725]/_0_  (.A(\inv_in[3725] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3726] ));
 sky130_fd_sc_hd__inv_2 \inv[3726]/_0_  (.A(\inv_in[3726] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3727] ));
 sky130_fd_sc_hd__inv_2 \inv[3727]/_0_  (.A(\inv_in[3727] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3728] ));
 sky130_fd_sc_hd__inv_2 \inv[3728]/_0_  (.A(\inv_in[3728] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3729] ));
 sky130_fd_sc_hd__inv_2 \inv[3729]/_0_  (.A(\inv_in[3729] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3730] ));
 sky130_fd_sc_hd__inv_2 \inv[372]/_0_  (.A(\inv_in[372] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[373] ));
 sky130_fd_sc_hd__inv_2 \inv[3730]/_0_  (.A(\inv_in[3730] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3731] ));
 sky130_fd_sc_hd__inv_2 \inv[3731]/_0_  (.A(\inv_in[3731] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3732] ));
 sky130_fd_sc_hd__inv_2 \inv[3732]/_0_  (.A(\inv_in[3732] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3733] ));
 sky130_fd_sc_hd__inv_2 \inv[3733]/_0_  (.A(\inv_in[3733] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3734] ));
 sky130_fd_sc_hd__inv_2 \inv[3734]/_0_  (.A(\inv_in[3734] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3735] ));
 sky130_fd_sc_hd__inv_2 \inv[3735]/_0_  (.A(\inv_in[3735] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3736] ));
 sky130_fd_sc_hd__inv_2 \inv[3736]/_0_  (.A(\inv_in[3736] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3737] ));
 sky130_fd_sc_hd__inv_2 \inv[3737]/_0_  (.A(\inv_in[3737] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3738] ));
 sky130_fd_sc_hd__inv_2 \inv[3738]/_0_  (.A(\inv_in[3738] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3739] ));
 sky130_fd_sc_hd__inv_2 \inv[3739]/_0_  (.A(\inv_in[3739] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3740] ));
 sky130_fd_sc_hd__inv_2 \inv[373]/_0_  (.A(\inv_in[373] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[374] ));
 sky130_fd_sc_hd__inv_2 \inv[3740]/_0_  (.A(\inv_in[3740] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3741] ));
 sky130_fd_sc_hd__inv_2 \inv[3741]/_0_  (.A(\inv_in[3741] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3742] ));
 sky130_fd_sc_hd__inv_2 \inv[3742]/_0_  (.A(\inv_in[3742] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3743] ));
 sky130_fd_sc_hd__inv_2 \inv[3743]/_0_  (.A(\inv_in[3743] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3744] ));
 sky130_fd_sc_hd__inv_2 \inv[3744]/_0_  (.A(\inv_in[3744] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3745] ));
 sky130_fd_sc_hd__inv_2 \inv[3745]/_0_  (.A(\inv_in[3745] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3746] ));
 sky130_fd_sc_hd__inv_2 \inv[3746]/_0_  (.A(\inv_in[3746] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3747] ));
 sky130_fd_sc_hd__inv_2 \inv[3747]/_0_  (.A(\inv_in[3747] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3748] ));
 sky130_fd_sc_hd__inv_2 \inv[3748]/_0_  (.A(\inv_in[3748] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3749] ));
 sky130_fd_sc_hd__inv_2 \inv[3749]/_0_  (.A(\inv_in[3749] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3750] ));
 sky130_fd_sc_hd__inv_2 \inv[374]/_0_  (.A(\inv_in[374] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[375] ));
 sky130_fd_sc_hd__inv_2 \inv[3750]/_0_  (.A(\inv_in[3750] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3751] ));
 sky130_fd_sc_hd__inv_2 \inv[3751]/_0_  (.A(\inv_in[3751] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3752] ));
 sky130_fd_sc_hd__inv_2 \inv[3752]/_0_  (.A(\inv_in[3752] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3753] ));
 sky130_fd_sc_hd__inv_2 \inv[3753]/_0_  (.A(\inv_in[3753] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3754] ));
 sky130_fd_sc_hd__inv_2 \inv[3754]/_0_  (.A(\inv_in[3754] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3755] ));
 sky130_fd_sc_hd__inv_2 \inv[3755]/_0_  (.A(\inv_in[3755] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3756] ));
 sky130_fd_sc_hd__inv_2 \inv[3756]/_0_  (.A(\inv_in[3756] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3757] ));
 sky130_fd_sc_hd__inv_2 \inv[3757]/_0_  (.A(\inv_in[3757] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3758] ));
 sky130_fd_sc_hd__inv_2 \inv[3758]/_0_  (.A(\inv_in[3758] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3759] ));
 sky130_fd_sc_hd__inv_2 \inv[3759]/_0_  (.A(\inv_in[3759] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3760] ));
 sky130_fd_sc_hd__inv_2 \inv[375]/_0_  (.A(\inv_in[375] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[376] ));
 sky130_fd_sc_hd__inv_2 \inv[3760]/_0_  (.A(\inv_in[3760] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3761] ));
 sky130_fd_sc_hd__inv_2 \inv[3761]/_0_  (.A(\inv_in[3761] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3762] ));
 sky130_fd_sc_hd__inv_2 \inv[3762]/_0_  (.A(\inv_in[3762] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3763] ));
 sky130_fd_sc_hd__inv_2 \inv[3763]/_0_  (.A(\inv_in[3763] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3764] ));
 sky130_fd_sc_hd__inv_2 \inv[3764]/_0_  (.A(\inv_in[3764] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3765] ));
 sky130_fd_sc_hd__inv_2 \inv[3765]/_0_  (.A(\inv_in[3765] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3766] ));
 sky130_fd_sc_hd__inv_2 \inv[3766]/_0_  (.A(\inv_in[3766] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3767] ));
 sky130_fd_sc_hd__inv_2 \inv[3767]/_0_  (.A(\inv_in[3767] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3768] ));
 sky130_fd_sc_hd__inv_2 \inv[3768]/_0_  (.A(\inv_in[3768] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3769] ));
 sky130_fd_sc_hd__inv_2 \inv[3769]/_0_  (.A(\inv_in[3769] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3770] ));
 sky130_fd_sc_hd__inv_2 \inv[376]/_0_  (.A(\inv_in[376] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[377] ));
 sky130_fd_sc_hd__inv_2 \inv[3770]/_0_  (.A(\inv_in[3770] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3771] ));
 sky130_fd_sc_hd__inv_2 \inv[3771]/_0_  (.A(\inv_in[3771] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3772] ));
 sky130_fd_sc_hd__inv_2 \inv[3772]/_0_  (.A(\inv_in[3772] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3773] ));
 sky130_fd_sc_hd__inv_2 \inv[3773]/_0_  (.A(\inv_in[3773] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3774] ));
 sky130_fd_sc_hd__inv_2 \inv[3774]/_0_  (.A(\inv_in[3774] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3775] ));
 sky130_fd_sc_hd__inv_2 \inv[3775]/_0_  (.A(\inv_in[3775] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3776] ));
 sky130_fd_sc_hd__inv_2 \inv[3776]/_0_  (.A(\inv_in[3776] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3777] ));
 sky130_fd_sc_hd__inv_2 \inv[3777]/_0_  (.A(\inv_in[3777] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3778] ));
 sky130_fd_sc_hd__inv_2 \inv[3778]/_0_  (.A(\inv_in[3778] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3779] ));
 sky130_fd_sc_hd__inv_2 \inv[3779]/_0_  (.A(\inv_in[3779] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3780] ));
 sky130_fd_sc_hd__inv_2 \inv[377]/_0_  (.A(\inv_in[377] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[378] ));
 sky130_fd_sc_hd__inv_2 \inv[3780]/_0_  (.A(\inv_in[3780] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3781] ));
 sky130_fd_sc_hd__inv_2 \inv[3781]/_0_  (.A(\inv_in[3781] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3782] ));
 sky130_fd_sc_hd__inv_2 \inv[3782]/_0_  (.A(\inv_in[3782] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3783] ));
 sky130_fd_sc_hd__inv_2 \inv[3783]/_0_  (.A(\inv_in[3783] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3784] ));
 sky130_fd_sc_hd__inv_2 \inv[3784]/_0_  (.A(\inv_in[3784] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3785] ));
 sky130_fd_sc_hd__inv_2 \inv[3785]/_0_  (.A(\inv_in[3785] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3786] ));
 sky130_fd_sc_hd__inv_2 \inv[3786]/_0_  (.A(\inv_in[3786] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3787] ));
 sky130_fd_sc_hd__inv_2 \inv[3787]/_0_  (.A(\inv_in[3787] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3788] ));
 sky130_fd_sc_hd__inv_2 \inv[3788]/_0_  (.A(\inv_in[3788] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3789] ));
 sky130_fd_sc_hd__inv_2 \inv[3789]/_0_  (.A(\inv_in[3789] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3790] ));
 sky130_fd_sc_hd__inv_2 \inv[378]/_0_  (.A(\inv_in[378] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[379] ));
 sky130_fd_sc_hd__inv_2 \inv[3790]/_0_  (.A(\inv_in[3790] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3791] ));
 sky130_fd_sc_hd__inv_2 \inv[3791]/_0_  (.A(\inv_in[3791] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3792] ));
 sky130_fd_sc_hd__inv_2 \inv[3792]/_0_  (.A(\inv_in[3792] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3793] ));
 sky130_fd_sc_hd__inv_2 \inv[3793]/_0_  (.A(\inv_in[3793] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3794] ));
 sky130_fd_sc_hd__inv_2 \inv[3794]/_0_  (.A(\inv_in[3794] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3795] ));
 sky130_fd_sc_hd__inv_2 \inv[3795]/_0_  (.A(\inv_in[3795] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3796] ));
 sky130_fd_sc_hd__inv_2 \inv[3796]/_0_  (.A(\inv_in[3796] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3797] ));
 sky130_fd_sc_hd__inv_2 \inv[3797]/_0_  (.A(\inv_in[3797] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3798] ));
 sky130_fd_sc_hd__inv_2 \inv[3798]/_0_  (.A(\inv_in[3798] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3799] ));
 sky130_fd_sc_hd__inv_2 \inv[3799]/_0_  (.A(\inv_in[3799] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3800] ));
 sky130_fd_sc_hd__inv_2 \inv[379]/_0_  (.A(\inv_in[379] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[380] ));
 sky130_fd_sc_hd__inv_2 \inv[37]/_0_  (.A(\inv_in[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[38] ));
 sky130_fd_sc_hd__inv_2 \inv[3800]/_0_  (.A(\inv_in[3800] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3801] ));
 sky130_fd_sc_hd__inv_2 \inv[3801]/_0_  (.A(\inv_in[3801] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3802] ));
 sky130_fd_sc_hd__inv_2 \inv[3802]/_0_  (.A(\inv_in[3802] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3803] ));
 sky130_fd_sc_hd__inv_2 \inv[3803]/_0_  (.A(\inv_in[3803] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3804] ));
 sky130_fd_sc_hd__inv_2 \inv[3804]/_0_  (.A(\inv_in[3804] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3805] ));
 sky130_fd_sc_hd__inv_2 \inv[3805]/_0_  (.A(\inv_in[3805] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3806] ));
 sky130_fd_sc_hd__inv_2 \inv[3806]/_0_  (.A(\inv_in[3806] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3807] ));
 sky130_fd_sc_hd__inv_2 \inv[3807]/_0_  (.A(\inv_in[3807] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3808] ));
 sky130_fd_sc_hd__inv_2 \inv[3808]/_0_  (.A(\inv_in[3808] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3809] ));
 sky130_fd_sc_hd__inv_2 \inv[3809]/_0_  (.A(\inv_in[3809] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3810] ));
 sky130_fd_sc_hd__inv_2 \inv[380]/_0_  (.A(\inv_in[380] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[381] ));
 sky130_fd_sc_hd__inv_2 \inv[3810]/_0_  (.A(\inv_in[3810] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3811] ));
 sky130_fd_sc_hd__inv_2 \inv[3811]/_0_  (.A(\inv_in[3811] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3812] ));
 sky130_fd_sc_hd__inv_2 \inv[3812]/_0_  (.A(\inv_in[3812] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3813] ));
 sky130_fd_sc_hd__inv_2 \inv[3813]/_0_  (.A(\inv_in[3813] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3814] ));
 sky130_fd_sc_hd__inv_2 \inv[3814]/_0_  (.A(\inv_in[3814] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3815] ));
 sky130_fd_sc_hd__inv_2 \inv[3815]/_0_  (.A(\inv_in[3815] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3816] ));
 sky130_fd_sc_hd__inv_2 \inv[3816]/_0_  (.A(\inv_in[3816] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3817] ));
 sky130_fd_sc_hd__inv_2 \inv[3817]/_0_  (.A(\inv_in[3817] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3818] ));
 sky130_fd_sc_hd__inv_2 \inv[3818]/_0_  (.A(\inv_in[3818] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3819] ));
 sky130_fd_sc_hd__inv_2 \inv[3819]/_0_  (.A(\inv_in[3819] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3820] ));
 sky130_fd_sc_hd__inv_2 \inv[381]/_0_  (.A(\inv_in[381] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[382] ));
 sky130_fd_sc_hd__inv_2 \inv[3820]/_0_  (.A(\inv_in[3820] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3821] ));
 sky130_fd_sc_hd__inv_2 \inv[3821]/_0_  (.A(\inv_in[3821] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3822] ));
 sky130_fd_sc_hd__inv_2 \inv[3822]/_0_  (.A(\inv_in[3822] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3823] ));
 sky130_fd_sc_hd__inv_2 \inv[3823]/_0_  (.A(\inv_in[3823] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3824] ));
 sky130_fd_sc_hd__inv_2 \inv[3824]/_0_  (.A(\inv_in[3824] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3825] ));
 sky130_fd_sc_hd__inv_2 \inv[3825]/_0_  (.A(\inv_in[3825] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3826] ));
 sky130_fd_sc_hd__inv_2 \inv[3826]/_0_  (.A(\inv_in[3826] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3827] ));
 sky130_fd_sc_hd__inv_2 \inv[3827]/_0_  (.A(\inv_in[3827] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3828] ));
 sky130_fd_sc_hd__inv_2 \inv[3828]/_0_  (.A(\inv_in[3828] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3829] ));
 sky130_fd_sc_hd__inv_2 \inv[3829]/_0_  (.A(\inv_in[3829] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3830] ));
 sky130_fd_sc_hd__inv_2 \inv[382]/_0_  (.A(\inv_in[382] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[383] ));
 sky130_fd_sc_hd__inv_2 \inv[3830]/_0_  (.A(\inv_in[3830] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3831] ));
 sky130_fd_sc_hd__inv_2 \inv[3831]/_0_  (.A(\inv_in[3831] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3832] ));
 sky130_fd_sc_hd__inv_2 \inv[3832]/_0_  (.A(\inv_in[3832] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3833] ));
 sky130_fd_sc_hd__inv_2 \inv[3833]/_0_  (.A(\inv_in[3833] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3834] ));
 sky130_fd_sc_hd__inv_2 \inv[3834]/_0_  (.A(\inv_in[3834] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3835] ));
 sky130_fd_sc_hd__inv_2 \inv[3835]/_0_  (.A(\inv_in[3835] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3836] ));
 sky130_fd_sc_hd__inv_2 \inv[3836]/_0_  (.A(\inv_in[3836] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3837] ));
 sky130_fd_sc_hd__inv_2 \inv[3837]/_0_  (.A(\inv_in[3837] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3838] ));
 sky130_fd_sc_hd__inv_2 \inv[3838]/_0_  (.A(\inv_in[3838] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3839] ));
 sky130_fd_sc_hd__inv_2 \inv[3839]/_0_  (.A(\inv_in[3839] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3840] ));
 sky130_fd_sc_hd__inv_2 \inv[383]/_0_  (.A(\inv_in[383] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[384] ));
 sky130_fd_sc_hd__inv_2 \inv[3840]/_0_  (.A(\inv_in[3840] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3841] ));
 sky130_fd_sc_hd__inv_2 \inv[3841]/_0_  (.A(\inv_in[3841] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3842] ));
 sky130_fd_sc_hd__inv_2 \inv[3842]/_0_  (.A(\inv_in[3842] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3843] ));
 sky130_fd_sc_hd__inv_2 \inv[3843]/_0_  (.A(\inv_in[3843] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3844] ));
 sky130_fd_sc_hd__inv_2 \inv[3844]/_0_  (.A(\inv_in[3844] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3845] ));
 sky130_fd_sc_hd__inv_2 \inv[3845]/_0_  (.A(\inv_in[3845] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3846] ));
 sky130_fd_sc_hd__inv_2 \inv[3846]/_0_  (.A(\inv_in[3846] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3847] ));
 sky130_fd_sc_hd__inv_2 \inv[3847]/_0_  (.A(\inv_in[3847] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3848] ));
 sky130_fd_sc_hd__inv_2 \inv[3848]/_0_  (.A(\inv_in[3848] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3849] ));
 sky130_fd_sc_hd__inv_2 \inv[3849]/_0_  (.A(\inv_in[3849] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3850] ));
 sky130_fd_sc_hd__inv_2 \inv[384]/_0_  (.A(\inv_in[384] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[385] ));
 sky130_fd_sc_hd__inv_2 \inv[3850]/_0_  (.A(\inv_in[3850] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3851] ));
 sky130_fd_sc_hd__inv_2 \inv[3851]/_0_  (.A(\inv_in[3851] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[3852] ));
 sky130_fd_sc_hd__inv_2 \inv[3852]/_0_  (.A(\inv_in[3852] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(uio_out[5]));
 sky130_fd_sc_hd__inv_2 \inv[385]/_0_  (.A(\inv_in[385] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[386] ));
 sky130_fd_sc_hd__inv_2 \inv[386]/_0_  (.A(\inv_in[386] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[387] ));
 sky130_fd_sc_hd__inv_2 \inv[387]/_0_  (.A(\inv_in[387] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[388] ));
 sky130_fd_sc_hd__inv_2 \inv[388]/_0_  (.A(\inv_in[388] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[389] ));
 sky130_fd_sc_hd__inv_2 \inv[389]/_0_  (.A(\inv_in[389] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[390] ));
 sky130_fd_sc_hd__inv_2 \inv[38]/_0_  (.A(\inv_in[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[39] ));
 sky130_fd_sc_hd__inv_2 \inv[390]/_0_  (.A(\inv_in[390] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[391] ));
 sky130_fd_sc_hd__inv_2 \inv[391]/_0_  (.A(\inv_in[391] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[392] ));
 sky130_fd_sc_hd__inv_2 \inv[392]/_0_  (.A(\inv_in[392] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[393] ));
 sky130_fd_sc_hd__inv_2 \inv[393]/_0_  (.A(\inv_in[393] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[394] ));
 sky130_fd_sc_hd__inv_2 \inv[394]/_0_  (.A(\inv_in[394] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[395] ));
 sky130_fd_sc_hd__inv_2 \inv[395]/_0_  (.A(\inv_in[395] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[396] ));
 sky130_fd_sc_hd__inv_2 \inv[396]/_0_  (.A(\inv_in[396] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[397] ));
 sky130_fd_sc_hd__inv_2 \inv[397]/_0_  (.A(\inv_in[397] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[398] ));
 sky130_fd_sc_hd__inv_2 \inv[398]/_0_  (.A(\inv_in[398] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[399] ));
 sky130_fd_sc_hd__inv_2 \inv[399]/_0_  (.A(\inv_in[399] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[400] ));
 sky130_fd_sc_hd__inv_2 \inv[39]/_0_  (.A(\inv_in[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[40] ));
 sky130_fd_sc_hd__inv_2 \inv[3]/_0_  (.A(\inv_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[4] ));
 sky130_fd_sc_hd__inv_2 \inv[400]/_0_  (.A(\inv_in[400] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[401] ));
 sky130_fd_sc_hd__inv_2 \inv[401]/_0_  (.A(\inv_in[401] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[402] ));
 sky130_fd_sc_hd__inv_2 \inv[402]/_0_  (.A(\inv_in[402] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[403] ));
 sky130_fd_sc_hd__inv_2 \inv[403]/_0_  (.A(\inv_in[403] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[404] ));
 sky130_fd_sc_hd__inv_2 \inv[404]/_0_  (.A(\inv_in[404] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[405] ));
 sky130_fd_sc_hd__inv_2 \inv[405]/_0_  (.A(\inv_in[405] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[406] ));
 sky130_fd_sc_hd__inv_2 \inv[406]/_0_  (.A(\inv_in[406] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[407] ));
 sky130_fd_sc_hd__inv_2 \inv[407]/_0_  (.A(\inv_in[407] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[408] ));
 sky130_fd_sc_hd__inv_2 \inv[408]/_0_  (.A(\inv_in[408] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[409] ));
 sky130_fd_sc_hd__inv_2 \inv[409]/_0_  (.A(\inv_in[409] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[410] ));
 sky130_fd_sc_hd__inv_2 \inv[40]/_0_  (.A(\inv_in[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[41] ));
 sky130_fd_sc_hd__inv_2 \inv[410]/_0_  (.A(\inv_in[410] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[411] ));
 sky130_fd_sc_hd__inv_2 \inv[411]/_0_  (.A(\inv_in[411] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[412] ));
 sky130_fd_sc_hd__inv_2 \inv[412]/_0_  (.A(\inv_in[412] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[413] ));
 sky130_fd_sc_hd__inv_2 \inv[413]/_0_  (.A(\inv_in[413] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[414] ));
 sky130_fd_sc_hd__inv_2 \inv[414]/_0_  (.A(\inv_in[414] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[415] ));
 sky130_fd_sc_hd__inv_2 \inv[415]/_0_  (.A(\inv_in[415] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[416] ));
 sky130_fd_sc_hd__inv_2 \inv[416]/_0_  (.A(\inv_in[416] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[417] ));
 sky130_fd_sc_hd__inv_2 \inv[417]/_0_  (.A(\inv_in[417] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[418] ));
 sky130_fd_sc_hd__inv_2 \inv[418]/_0_  (.A(\inv_in[418] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[419] ));
 sky130_fd_sc_hd__inv_2 \inv[419]/_0_  (.A(\inv_in[419] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[420] ));
 sky130_fd_sc_hd__inv_2 \inv[41]/_0_  (.A(\inv_in[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[42] ));
 sky130_fd_sc_hd__inv_2 \inv[420]/_0_  (.A(\inv_in[420] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[421] ));
 sky130_fd_sc_hd__inv_2 \inv[421]/_0_  (.A(\inv_in[421] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[422] ));
 sky130_fd_sc_hd__inv_2 \inv[422]/_0_  (.A(\inv_in[422] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[423] ));
 sky130_fd_sc_hd__inv_2 \inv[423]/_0_  (.A(\inv_in[423] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[424] ));
 sky130_fd_sc_hd__inv_2 \inv[424]/_0_  (.A(\inv_in[424] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[425] ));
 sky130_fd_sc_hd__inv_2 \inv[425]/_0_  (.A(\inv_in[425] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[426] ));
 sky130_fd_sc_hd__inv_2 \inv[426]/_0_  (.A(\inv_in[426] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[427] ));
 sky130_fd_sc_hd__inv_2 \inv[427]/_0_  (.A(\inv_in[427] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[428] ));
 sky130_fd_sc_hd__inv_2 \inv[428]/_0_  (.A(\inv_in[428] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[429] ));
 sky130_fd_sc_hd__inv_2 \inv[429]/_0_  (.A(\inv_in[429] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[430] ));
 sky130_fd_sc_hd__inv_2 \inv[42]/_0_  (.A(\inv_in[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[43] ));
 sky130_fd_sc_hd__inv_2 \inv[430]/_0_  (.A(\inv_in[430] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[431] ));
 sky130_fd_sc_hd__inv_2 \inv[431]/_0_  (.A(\inv_in[431] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[432] ));
 sky130_fd_sc_hd__inv_2 \inv[432]/_0_  (.A(\inv_in[432] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[433] ));
 sky130_fd_sc_hd__inv_2 \inv[433]/_0_  (.A(\inv_in[433] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[434] ));
 sky130_fd_sc_hd__inv_2 \inv[434]/_0_  (.A(\inv_in[434] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[435] ));
 sky130_fd_sc_hd__inv_2 \inv[435]/_0_  (.A(\inv_in[435] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[436] ));
 sky130_fd_sc_hd__inv_2 \inv[436]/_0_  (.A(\inv_in[436] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[437] ));
 sky130_fd_sc_hd__inv_2 \inv[437]/_0_  (.A(\inv_in[437] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[438] ));
 sky130_fd_sc_hd__inv_2 \inv[438]/_0_  (.A(\inv_in[438] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[439] ));
 sky130_fd_sc_hd__inv_2 \inv[439]/_0_  (.A(\inv_in[439] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[440] ));
 sky130_fd_sc_hd__inv_2 \inv[43]/_0_  (.A(\inv_in[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[44] ));
 sky130_fd_sc_hd__inv_2 \inv[440]/_0_  (.A(\inv_in[440] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[441] ));
 sky130_fd_sc_hd__inv_2 \inv[441]/_0_  (.A(\inv_in[441] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[442] ));
 sky130_fd_sc_hd__inv_2 \inv[442]/_0_  (.A(\inv_in[442] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[443] ));
 sky130_fd_sc_hd__inv_2 \inv[443]/_0_  (.A(\inv_in[443] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[444] ));
 sky130_fd_sc_hd__inv_2 \inv[444]/_0_  (.A(\inv_in[444] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[445] ));
 sky130_fd_sc_hd__inv_2 \inv[445]/_0_  (.A(\inv_in[445] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[446] ));
 sky130_fd_sc_hd__inv_2 \inv[446]/_0_  (.A(\inv_in[446] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[447] ));
 sky130_fd_sc_hd__inv_2 \inv[447]/_0_  (.A(\inv_in[447] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[448] ));
 sky130_fd_sc_hd__inv_2 \inv[448]/_0_  (.A(\inv_in[448] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[449] ));
 sky130_fd_sc_hd__inv_2 \inv[449]/_0_  (.A(\inv_in[449] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[450] ));
 sky130_fd_sc_hd__inv_2 \inv[44]/_0_  (.A(\inv_in[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[45] ));
 sky130_fd_sc_hd__inv_2 \inv[450]/_0_  (.A(\inv_in[450] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[451] ));
 sky130_fd_sc_hd__inv_2 \inv[451]/_0_  (.A(\inv_in[451] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[452] ));
 sky130_fd_sc_hd__inv_2 \inv[452]/_0_  (.A(\inv_in[452] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[453] ));
 sky130_fd_sc_hd__inv_2 \inv[453]/_0_  (.A(\inv_in[453] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[454] ));
 sky130_fd_sc_hd__inv_2 \inv[454]/_0_  (.A(\inv_in[454] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[455] ));
 sky130_fd_sc_hd__inv_2 \inv[455]/_0_  (.A(\inv_in[455] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[456] ));
 sky130_fd_sc_hd__inv_2 \inv[456]/_0_  (.A(\inv_in[456] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[457] ));
 sky130_fd_sc_hd__inv_2 \inv[457]/_0_  (.A(\inv_in[457] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[458] ));
 sky130_fd_sc_hd__inv_2 \inv[458]/_0_  (.A(\inv_in[458] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[459] ));
 sky130_fd_sc_hd__inv_2 \inv[459]/_0_  (.A(\inv_in[459] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[460] ));
 sky130_fd_sc_hd__inv_2 \inv[45]/_0_  (.A(\inv_in[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[46] ));
 sky130_fd_sc_hd__inv_2 \inv[460]/_0_  (.A(\inv_in[460] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[461] ));
 sky130_fd_sc_hd__inv_2 \inv[461]/_0_  (.A(\inv_in[461] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[462] ));
 sky130_fd_sc_hd__inv_2 \inv[462]/_0_  (.A(\inv_in[462] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[463] ));
 sky130_fd_sc_hd__inv_2 \inv[463]/_0_  (.A(\inv_in[463] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[464] ));
 sky130_fd_sc_hd__inv_2 \inv[464]/_0_  (.A(\inv_in[464] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[465] ));
 sky130_fd_sc_hd__inv_2 \inv[465]/_0_  (.A(\inv_in[465] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[466] ));
 sky130_fd_sc_hd__inv_2 \inv[466]/_0_  (.A(\inv_in[466] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[467] ));
 sky130_fd_sc_hd__inv_2 \inv[467]/_0_  (.A(\inv_in[467] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[468] ));
 sky130_fd_sc_hd__inv_2 \inv[468]/_0_  (.A(\inv_in[468] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[469] ));
 sky130_fd_sc_hd__inv_2 \inv[469]/_0_  (.A(\inv_in[469] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[470] ));
 sky130_fd_sc_hd__inv_2 \inv[46]/_0_  (.A(\inv_in[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[47] ));
 sky130_fd_sc_hd__inv_2 \inv[470]/_0_  (.A(\inv_in[470] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[471] ));
 sky130_fd_sc_hd__inv_2 \inv[471]/_0_  (.A(\inv_in[471] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[472] ));
 sky130_fd_sc_hd__inv_2 \inv[472]/_0_  (.A(\inv_in[472] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[473] ));
 sky130_fd_sc_hd__inv_2 \inv[473]/_0_  (.A(\inv_in[473] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[474] ));
 sky130_fd_sc_hd__inv_2 \inv[474]/_0_  (.A(\inv_in[474] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[475] ));
 sky130_fd_sc_hd__inv_2 \inv[475]/_0_  (.A(\inv_in[475] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[476] ));
 sky130_fd_sc_hd__inv_2 \inv[476]/_0_  (.A(\inv_in[476] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[477] ));
 sky130_fd_sc_hd__inv_2 \inv[477]/_0_  (.A(\inv_in[477] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[478] ));
 sky130_fd_sc_hd__inv_2 \inv[478]/_0_  (.A(\inv_in[478] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[479] ));
 sky130_fd_sc_hd__inv_2 \inv[479]/_0_  (.A(\inv_in[479] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[480] ));
 sky130_fd_sc_hd__inv_2 \inv[47]/_0_  (.A(\inv_in[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[48] ));
 sky130_fd_sc_hd__inv_2 \inv[480]/_0_  (.A(\inv_in[480] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[481] ));
 sky130_fd_sc_hd__inv_2 \inv[481]/_0_  (.A(\inv_in[481] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[482] ));
 sky130_fd_sc_hd__inv_2 \inv[482]/_0_  (.A(\inv_in[482] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[483] ));
 sky130_fd_sc_hd__inv_2 \inv[483]/_0_  (.A(\inv_in[483] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[484] ));
 sky130_fd_sc_hd__inv_2 \inv[484]/_0_  (.A(\inv_in[484] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[485] ));
 sky130_fd_sc_hd__inv_2 \inv[485]/_0_  (.A(\inv_in[485] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[486] ));
 sky130_fd_sc_hd__inv_2 \inv[486]/_0_  (.A(\inv_in[486] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[487] ));
 sky130_fd_sc_hd__inv_2 \inv[487]/_0_  (.A(\inv_in[487] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[488] ));
 sky130_fd_sc_hd__inv_2 \inv[488]/_0_  (.A(\inv_in[488] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[489] ));
 sky130_fd_sc_hd__inv_2 \inv[489]/_0_  (.A(\inv_in[489] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[490] ));
 sky130_fd_sc_hd__inv_2 \inv[48]/_0_  (.A(\inv_in[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[49] ));
 sky130_fd_sc_hd__inv_2 \inv[490]/_0_  (.A(\inv_in[490] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[491] ));
 sky130_fd_sc_hd__inv_2 \inv[491]/_0_  (.A(\inv_in[491] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[492] ));
 sky130_fd_sc_hd__inv_2 \inv[492]/_0_  (.A(\inv_in[492] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[493] ));
 sky130_fd_sc_hd__inv_2 \inv[493]/_0_  (.A(\inv_in[493] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[494] ));
 sky130_fd_sc_hd__inv_2 \inv[494]/_0_  (.A(\inv_in[494] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[495] ));
 sky130_fd_sc_hd__inv_2 \inv[495]/_0_  (.A(\inv_in[495] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[496] ));
 sky130_fd_sc_hd__inv_2 \inv[496]/_0_  (.A(\inv_in[496] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[497] ));
 sky130_fd_sc_hd__inv_2 \inv[497]/_0_  (.A(\inv_in[497] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[498] ));
 sky130_fd_sc_hd__inv_2 \inv[498]/_0_  (.A(\inv_in[498] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[499] ));
 sky130_fd_sc_hd__inv_2 \inv[499]/_0_  (.A(\inv_in[499] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[500] ));
 sky130_fd_sc_hd__inv_2 \inv[49]/_0_  (.A(\inv_in[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[50] ));
 sky130_fd_sc_hd__inv_2 \inv[4]/_0_  (.A(\inv_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[5] ));
 sky130_fd_sc_hd__inv_2 \inv[500]/_0_  (.A(\inv_in[500] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[501] ));
 sky130_fd_sc_hd__inv_2 \inv[501]/_0_  (.A(\inv_in[501] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[502] ));
 sky130_fd_sc_hd__inv_2 \inv[502]/_0_  (.A(\inv_in[502] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[503] ));
 sky130_fd_sc_hd__inv_2 \inv[503]/_0_  (.A(\inv_in[503] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[504] ));
 sky130_fd_sc_hd__inv_2 \inv[504]/_0_  (.A(\inv_in[504] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[505] ));
 sky130_fd_sc_hd__inv_2 \inv[505]/_0_  (.A(\inv_in[505] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[506] ));
 sky130_fd_sc_hd__inv_2 \inv[506]/_0_  (.A(\inv_in[506] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[507] ));
 sky130_fd_sc_hd__inv_2 \inv[507]/_0_  (.A(\inv_in[507] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[508] ));
 sky130_fd_sc_hd__inv_2 \inv[508]/_0_  (.A(\inv_in[508] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[509] ));
 sky130_fd_sc_hd__inv_2 \inv[509]/_0_  (.A(\inv_in[509] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[510] ));
 sky130_fd_sc_hd__inv_2 \inv[50]/_0_  (.A(\inv_in[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[51] ));
 sky130_fd_sc_hd__inv_2 \inv[510]/_0_  (.A(\inv_in[510] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[511] ));
 sky130_fd_sc_hd__inv_2 \inv[511]/_0_  (.A(\inv_in[511] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[512] ));
 sky130_fd_sc_hd__inv_2 \inv[512]/_0_  (.A(\inv_in[512] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[513] ));
 sky130_fd_sc_hd__inv_2 \inv[513]/_0_  (.A(\inv_in[513] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[514] ));
 sky130_fd_sc_hd__inv_2 \inv[514]/_0_  (.A(\inv_in[514] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[515] ));
 sky130_fd_sc_hd__inv_2 \inv[515]/_0_  (.A(\inv_in[515] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[516] ));
 sky130_fd_sc_hd__inv_2 \inv[516]/_0_  (.A(\inv_in[516] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[517] ));
 sky130_fd_sc_hd__inv_2 \inv[517]/_0_  (.A(\inv_in[517] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[518] ));
 sky130_fd_sc_hd__inv_2 \inv[518]/_0_  (.A(\inv_in[518] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[519] ));
 sky130_fd_sc_hd__inv_2 \inv[519]/_0_  (.A(\inv_in[519] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[520] ));
 sky130_fd_sc_hd__inv_2 \inv[51]/_0_  (.A(\inv_in[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[52] ));
 sky130_fd_sc_hd__inv_2 \inv[520]/_0_  (.A(\inv_in[520] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[521] ));
 sky130_fd_sc_hd__inv_2 \inv[521]/_0_  (.A(\inv_in[521] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[522] ));
 sky130_fd_sc_hd__inv_2 \inv[522]/_0_  (.A(\inv_in[522] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[523] ));
 sky130_fd_sc_hd__inv_2 \inv[523]/_0_  (.A(\inv_in[523] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[524] ));
 sky130_fd_sc_hd__inv_2 \inv[524]/_0_  (.A(\inv_in[524] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[525] ));
 sky130_fd_sc_hd__inv_2 \inv[525]/_0_  (.A(\inv_in[525] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[526] ));
 sky130_fd_sc_hd__inv_2 \inv[526]/_0_  (.A(\inv_in[526] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[527] ));
 sky130_fd_sc_hd__inv_2 \inv[527]/_0_  (.A(\inv_in[527] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[528] ));
 sky130_fd_sc_hd__inv_2 \inv[528]/_0_  (.A(\inv_in[528] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[529] ));
 sky130_fd_sc_hd__inv_2 \inv[529]/_0_  (.A(\inv_in[529] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[530] ));
 sky130_fd_sc_hd__inv_2 \inv[52]/_0_  (.A(\inv_in[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[53] ));
 sky130_fd_sc_hd__inv_2 \inv[530]/_0_  (.A(\inv_in[530] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[531] ));
 sky130_fd_sc_hd__inv_2 \inv[531]/_0_  (.A(\inv_in[531] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[532] ));
 sky130_fd_sc_hd__inv_2 \inv[532]/_0_  (.A(\inv_in[532] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[533] ));
 sky130_fd_sc_hd__inv_2 \inv[533]/_0_  (.A(\inv_in[533] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[534] ));
 sky130_fd_sc_hd__inv_2 \inv[534]/_0_  (.A(\inv_in[534] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[535] ));
 sky130_fd_sc_hd__inv_2 \inv[535]/_0_  (.A(\inv_in[535] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[536] ));
 sky130_fd_sc_hd__inv_2 \inv[536]/_0_  (.A(\inv_in[536] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[537] ));
 sky130_fd_sc_hd__inv_2 \inv[537]/_0_  (.A(\inv_in[537] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[538] ));
 sky130_fd_sc_hd__inv_2 \inv[538]/_0_  (.A(\inv_in[538] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[539] ));
 sky130_fd_sc_hd__inv_2 \inv[539]/_0_  (.A(\inv_in[539] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[540] ));
 sky130_fd_sc_hd__inv_2 \inv[53]/_0_  (.A(\inv_in[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[54] ));
 sky130_fd_sc_hd__inv_2 \inv[540]/_0_  (.A(\inv_in[540] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[541] ));
 sky130_fd_sc_hd__inv_2 \inv[541]/_0_  (.A(\inv_in[541] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[542] ));
 sky130_fd_sc_hd__inv_2 \inv[542]/_0_  (.A(\inv_in[542] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[543] ));
 sky130_fd_sc_hd__inv_2 \inv[543]/_0_  (.A(\inv_in[543] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[544] ));
 sky130_fd_sc_hd__inv_2 \inv[544]/_0_  (.A(\inv_in[544] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[545] ));
 sky130_fd_sc_hd__inv_2 \inv[545]/_0_  (.A(\inv_in[545] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[546] ));
 sky130_fd_sc_hd__inv_2 \inv[546]/_0_  (.A(\inv_in[546] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[547] ));
 sky130_fd_sc_hd__inv_2 \inv[547]/_0_  (.A(\inv_in[547] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[548] ));
 sky130_fd_sc_hd__inv_2 \inv[548]/_0_  (.A(\inv_in[548] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[549] ));
 sky130_fd_sc_hd__inv_2 \inv[549]/_0_  (.A(\inv_in[549] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[550] ));
 sky130_fd_sc_hd__inv_2 \inv[54]/_0_  (.A(\inv_in[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[55] ));
 sky130_fd_sc_hd__inv_2 \inv[550]/_0_  (.A(\inv_in[550] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[551] ));
 sky130_fd_sc_hd__inv_2 \inv[551]/_0_  (.A(\inv_in[551] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[552] ));
 sky130_fd_sc_hd__inv_2 \inv[552]/_0_  (.A(\inv_in[552] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[553] ));
 sky130_fd_sc_hd__inv_2 \inv[553]/_0_  (.A(\inv_in[553] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[554] ));
 sky130_fd_sc_hd__inv_2 \inv[554]/_0_  (.A(\inv_in[554] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[555] ));
 sky130_fd_sc_hd__inv_2 \inv[555]/_0_  (.A(\inv_in[555] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[556] ));
 sky130_fd_sc_hd__inv_2 \inv[556]/_0_  (.A(\inv_in[556] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[557] ));
 sky130_fd_sc_hd__inv_2 \inv[557]/_0_  (.A(\inv_in[557] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[558] ));
 sky130_fd_sc_hd__inv_2 \inv[558]/_0_  (.A(\inv_in[558] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[559] ));
 sky130_fd_sc_hd__inv_2 \inv[559]/_0_  (.A(\inv_in[559] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[560] ));
 sky130_fd_sc_hd__inv_2 \inv[55]/_0_  (.A(\inv_in[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[56] ));
 sky130_fd_sc_hd__inv_2 \inv[560]/_0_  (.A(\inv_in[560] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[561] ));
 sky130_fd_sc_hd__inv_2 \inv[561]/_0_  (.A(\inv_in[561] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[562] ));
 sky130_fd_sc_hd__inv_2 \inv[562]/_0_  (.A(\inv_in[562] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[563] ));
 sky130_fd_sc_hd__inv_2 \inv[563]/_0_  (.A(\inv_in[563] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[564] ));
 sky130_fd_sc_hd__inv_2 \inv[564]/_0_  (.A(\inv_in[564] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[565] ));
 sky130_fd_sc_hd__inv_2 \inv[565]/_0_  (.A(\inv_in[565] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[566] ));
 sky130_fd_sc_hd__inv_2 \inv[566]/_0_  (.A(\inv_in[566] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[567] ));
 sky130_fd_sc_hd__inv_2 \inv[567]/_0_  (.A(\inv_in[567] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[568] ));
 sky130_fd_sc_hd__inv_2 \inv[568]/_0_  (.A(\inv_in[568] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[569] ));
 sky130_fd_sc_hd__inv_2 \inv[569]/_0_  (.A(\inv_in[569] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[570] ));
 sky130_fd_sc_hd__inv_2 \inv[56]/_0_  (.A(\inv_in[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[57] ));
 sky130_fd_sc_hd__inv_2 \inv[570]/_0_  (.A(\inv_in[570] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[571] ));
 sky130_fd_sc_hd__inv_2 \inv[571]/_0_  (.A(\inv_in[571] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[572] ));
 sky130_fd_sc_hd__inv_2 \inv[572]/_0_  (.A(\inv_in[572] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[573] ));
 sky130_fd_sc_hd__inv_2 \inv[573]/_0_  (.A(\inv_in[573] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[574] ));
 sky130_fd_sc_hd__inv_2 \inv[574]/_0_  (.A(\inv_in[574] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[575] ));
 sky130_fd_sc_hd__inv_2 \inv[575]/_0_  (.A(\inv_in[575] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[576] ));
 sky130_fd_sc_hd__inv_2 \inv[576]/_0_  (.A(\inv_in[576] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[577] ));
 sky130_fd_sc_hd__inv_2 \inv[577]/_0_  (.A(\inv_in[577] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[578] ));
 sky130_fd_sc_hd__inv_2 \inv[578]/_0_  (.A(\inv_in[578] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[579] ));
 sky130_fd_sc_hd__inv_2 \inv[579]/_0_  (.A(\inv_in[579] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[580] ));
 sky130_fd_sc_hd__inv_2 \inv[57]/_0_  (.A(\inv_in[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[58] ));
 sky130_fd_sc_hd__inv_2 \inv[580]/_0_  (.A(\inv_in[580] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[581] ));
 sky130_fd_sc_hd__inv_2 \inv[581]/_0_  (.A(\inv_in[581] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[582] ));
 sky130_fd_sc_hd__inv_2 \inv[582]/_0_  (.A(\inv_in[582] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[583] ));
 sky130_fd_sc_hd__inv_2 \inv[583]/_0_  (.A(\inv_in[583] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[584] ));
 sky130_fd_sc_hd__inv_2 \inv[584]/_0_  (.A(\inv_in[584] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[585] ));
 sky130_fd_sc_hd__inv_2 \inv[585]/_0_  (.A(\inv_in[585] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[586] ));
 sky130_fd_sc_hd__inv_2 \inv[586]/_0_  (.A(\inv_in[586] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[587] ));
 sky130_fd_sc_hd__inv_2 \inv[587]/_0_  (.A(\inv_in[587] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[588] ));
 sky130_fd_sc_hd__inv_2 \inv[588]/_0_  (.A(\inv_in[588] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[589] ));
 sky130_fd_sc_hd__inv_2 \inv[589]/_0_  (.A(\inv_in[589] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[590] ));
 sky130_fd_sc_hd__inv_2 \inv[58]/_0_  (.A(\inv_in[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[59] ));
 sky130_fd_sc_hd__inv_2 \inv[590]/_0_  (.A(\inv_in[590] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[591] ));
 sky130_fd_sc_hd__inv_2 \inv[591]/_0_  (.A(\inv_in[591] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[592] ));
 sky130_fd_sc_hd__inv_2 \inv[592]/_0_  (.A(\inv_in[592] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[593] ));
 sky130_fd_sc_hd__inv_2 \inv[593]/_0_  (.A(\inv_in[593] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[594] ));
 sky130_fd_sc_hd__inv_2 \inv[594]/_0_  (.A(\inv_in[594] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[595] ));
 sky130_fd_sc_hd__inv_2 \inv[595]/_0_  (.A(\inv_in[595] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[596] ));
 sky130_fd_sc_hd__inv_2 \inv[596]/_0_  (.A(\inv_in[596] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[597] ));
 sky130_fd_sc_hd__inv_2 \inv[597]/_0_  (.A(\inv_in[597] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[598] ));
 sky130_fd_sc_hd__inv_2 \inv[598]/_0_  (.A(\inv_in[598] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[599] ));
 sky130_fd_sc_hd__inv_2 \inv[599]/_0_  (.A(\inv_in[599] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[600] ));
 sky130_fd_sc_hd__inv_2 \inv[59]/_0_  (.A(\inv_in[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[60] ));
 sky130_fd_sc_hd__inv_2 \inv[5]/_0_  (.A(\inv_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[6] ));
 sky130_fd_sc_hd__inv_2 \inv[600]/_0_  (.A(\inv_in[600] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[601] ));
 sky130_fd_sc_hd__inv_2 \inv[601]/_0_  (.A(\inv_in[601] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[602] ));
 sky130_fd_sc_hd__inv_2 \inv[602]/_0_  (.A(\inv_in[602] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[603] ));
 sky130_fd_sc_hd__inv_2 \inv[603]/_0_  (.A(\inv_in[603] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[604] ));
 sky130_fd_sc_hd__inv_2 \inv[604]/_0_  (.A(\inv_in[604] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[605] ));
 sky130_fd_sc_hd__inv_2 \inv[605]/_0_  (.A(\inv_in[605] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[606] ));
 sky130_fd_sc_hd__inv_2 \inv[606]/_0_  (.A(\inv_in[606] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[607] ));
 sky130_fd_sc_hd__inv_2 \inv[607]/_0_  (.A(\inv_in[607] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[608] ));
 sky130_fd_sc_hd__inv_2 \inv[608]/_0_  (.A(\inv_in[608] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[609] ));
 sky130_fd_sc_hd__inv_2 \inv[609]/_0_  (.A(\inv_in[609] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[610] ));
 sky130_fd_sc_hd__inv_2 \inv[60]/_0_  (.A(\inv_in[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[61] ));
 sky130_fd_sc_hd__inv_2 \inv[610]/_0_  (.A(\inv_in[610] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[611] ));
 sky130_fd_sc_hd__inv_2 \inv[611]/_0_  (.A(\inv_in[611] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[612] ));
 sky130_fd_sc_hd__inv_2 \inv[612]/_0_  (.A(\inv_in[612] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[613] ));
 sky130_fd_sc_hd__inv_2 \inv[613]/_0_  (.A(\inv_in[613] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[614] ));
 sky130_fd_sc_hd__inv_2 \inv[614]/_0_  (.A(\inv_in[614] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[615] ));
 sky130_fd_sc_hd__inv_2 \inv[615]/_0_  (.A(\inv_in[615] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[616] ));
 sky130_fd_sc_hd__inv_2 \inv[616]/_0_  (.A(\inv_in[616] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[617] ));
 sky130_fd_sc_hd__inv_2 \inv[617]/_0_  (.A(\inv_in[617] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[618] ));
 sky130_fd_sc_hd__inv_2 \inv[618]/_0_  (.A(\inv_in[618] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[619] ));
 sky130_fd_sc_hd__inv_2 \inv[619]/_0_  (.A(\inv_in[619] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[620] ));
 sky130_fd_sc_hd__inv_2 \inv[61]/_0_  (.A(\inv_in[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[62] ));
 sky130_fd_sc_hd__inv_2 \inv[620]/_0_  (.A(\inv_in[620] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[621] ));
 sky130_fd_sc_hd__inv_2 \inv[621]/_0_  (.A(\inv_in[621] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[622] ));
 sky130_fd_sc_hd__inv_2 \inv[622]/_0_  (.A(\inv_in[622] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[623] ));
 sky130_fd_sc_hd__inv_2 \inv[623]/_0_  (.A(\inv_in[623] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[624] ));
 sky130_fd_sc_hd__inv_2 \inv[624]/_0_  (.A(\inv_in[624] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[625] ));
 sky130_fd_sc_hd__inv_2 \inv[625]/_0_  (.A(\inv_in[625] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[626] ));
 sky130_fd_sc_hd__inv_2 \inv[626]/_0_  (.A(\inv_in[626] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[627] ));
 sky130_fd_sc_hd__inv_2 \inv[627]/_0_  (.A(\inv_in[627] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[628] ));
 sky130_fd_sc_hd__inv_2 \inv[628]/_0_  (.A(\inv_in[628] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[629] ));
 sky130_fd_sc_hd__inv_2 \inv[629]/_0_  (.A(\inv_in[629] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[630] ));
 sky130_fd_sc_hd__inv_2 \inv[62]/_0_  (.A(\inv_in[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[63] ));
 sky130_fd_sc_hd__inv_2 \inv[630]/_0_  (.A(\inv_in[630] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[631] ));
 sky130_fd_sc_hd__inv_2 \inv[631]/_0_  (.A(\inv_in[631] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[632] ));
 sky130_fd_sc_hd__inv_2 \inv[632]/_0_  (.A(\inv_in[632] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[633] ));
 sky130_fd_sc_hd__inv_2 \inv[633]/_0_  (.A(\inv_in[633] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[634] ));
 sky130_fd_sc_hd__inv_2 \inv[634]/_0_  (.A(\inv_in[634] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[635] ));
 sky130_fd_sc_hd__inv_2 \inv[635]/_0_  (.A(\inv_in[635] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[636] ));
 sky130_fd_sc_hd__inv_2 \inv[636]/_0_  (.A(\inv_in[636] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[637] ));
 sky130_fd_sc_hd__inv_2 \inv[637]/_0_  (.A(\inv_in[637] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[638] ));
 sky130_fd_sc_hd__inv_2 \inv[638]/_0_  (.A(\inv_in[638] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[639] ));
 sky130_fd_sc_hd__inv_2 \inv[639]/_0_  (.A(\inv_in[639] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[640] ));
 sky130_fd_sc_hd__inv_2 \inv[63]/_0_  (.A(\inv_in[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[64] ));
 sky130_fd_sc_hd__inv_2 \inv[640]/_0_  (.A(\inv_in[640] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[641] ));
 sky130_fd_sc_hd__inv_2 \inv[641]/_0_  (.A(\inv_in[641] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[642] ));
 sky130_fd_sc_hd__inv_2 \inv[642]/_0_  (.A(\inv_in[642] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[643] ));
 sky130_fd_sc_hd__inv_2 \inv[643]/_0_  (.A(\inv_in[643] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[644] ));
 sky130_fd_sc_hd__inv_2 \inv[644]/_0_  (.A(\inv_in[644] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[645] ));
 sky130_fd_sc_hd__inv_2 \inv[645]/_0_  (.A(\inv_in[645] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[646] ));
 sky130_fd_sc_hd__inv_2 \inv[646]/_0_  (.A(\inv_in[646] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[647] ));
 sky130_fd_sc_hd__inv_2 \inv[647]/_0_  (.A(\inv_in[647] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[648] ));
 sky130_fd_sc_hd__inv_2 \inv[648]/_0_  (.A(\inv_in[648] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[649] ));
 sky130_fd_sc_hd__inv_2 \inv[649]/_0_  (.A(\inv_in[649] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[650] ));
 sky130_fd_sc_hd__inv_2 \inv[64]/_0_  (.A(\inv_in[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[65] ));
 sky130_fd_sc_hd__inv_2 \inv[650]/_0_  (.A(\inv_in[650] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[651] ));
 sky130_fd_sc_hd__inv_2 \inv[651]/_0_  (.A(\inv_in[651] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[652] ));
 sky130_fd_sc_hd__inv_2 \inv[652]/_0_  (.A(\inv_in[652] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[653] ));
 sky130_fd_sc_hd__inv_2 \inv[653]/_0_  (.A(\inv_in[653] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[654] ));
 sky130_fd_sc_hd__inv_2 \inv[654]/_0_  (.A(\inv_in[654] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[655] ));
 sky130_fd_sc_hd__inv_2 \inv[655]/_0_  (.A(\inv_in[655] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[656] ));
 sky130_fd_sc_hd__inv_2 \inv[656]/_0_  (.A(\inv_in[656] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[657] ));
 sky130_fd_sc_hd__inv_2 \inv[657]/_0_  (.A(\inv_in[657] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[658] ));
 sky130_fd_sc_hd__inv_2 \inv[658]/_0_  (.A(\inv_in[658] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[659] ));
 sky130_fd_sc_hd__inv_2 \inv[659]/_0_  (.A(\inv_in[659] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[660] ));
 sky130_fd_sc_hd__inv_2 \inv[65]/_0_  (.A(\inv_in[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[66] ));
 sky130_fd_sc_hd__inv_2 \inv[660]/_0_  (.A(\inv_in[660] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[661] ));
 sky130_fd_sc_hd__inv_2 \inv[661]/_0_  (.A(\inv_in[661] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[662] ));
 sky130_fd_sc_hd__inv_2 \inv[662]/_0_  (.A(\inv_in[662] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[663] ));
 sky130_fd_sc_hd__inv_2 \inv[663]/_0_  (.A(\inv_in[663] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[664] ));
 sky130_fd_sc_hd__inv_2 \inv[664]/_0_  (.A(\inv_in[664] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[665] ));
 sky130_fd_sc_hd__inv_2 \inv[665]/_0_  (.A(\inv_in[665] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[666] ));
 sky130_fd_sc_hd__inv_2 \inv[666]/_0_  (.A(\inv_in[666] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[667] ));
 sky130_fd_sc_hd__inv_2 \inv[667]/_0_  (.A(\inv_in[667] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[668] ));
 sky130_fd_sc_hd__inv_2 \inv[668]/_0_  (.A(\inv_in[668] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[669] ));
 sky130_fd_sc_hd__inv_2 \inv[669]/_0_  (.A(\inv_in[669] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[670] ));
 sky130_fd_sc_hd__inv_2 \inv[66]/_0_  (.A(\inv_in[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[67] ));
 sky130_fd_sc_hd__inv_2 \inv[670]/_0_  (.A(\inv_in[670] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[671] ));
 sky130_fd_sc_hd__inv_2 \inv[671]/_0_  (.A(\inv_in[671] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[672] ));
 sky130_fd_sc_hd__inv_2 \inv[672]/_0_  (.A(\inv_in[672] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[673] ));
 sky130_fd_sc_hd__inv_2 \inv[673]/_0_  (.A(\inv_in[673] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[674] ));
 sky130_fd_sc_hd__inv_2 \inv[674]/_0_  (.A(\inv_in[674] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[675] ));
 sky130_fd_sc_hd__inv_2 \inv[675]/_0_  (.A(\inv_in[675] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[676] ));
 sky130_fd_sc_hd__inv_2 \inv[676]/_0_  (.A(\inv_in[676] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[677] ));
 sky130_fd_sc_hd__inv_2 \inv[677]/_0_  (.A(\inv_in[677] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[678] ));
 sky130_fd_sc_hd__inv_2 \inv[678]/_0_  (.A(\inv_in[678] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[679] ));
 sky130_fd_sc_hd__inv_2 \inv[679]/_0_  (.A(\inv_in[679] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[680] ));
 sky130_fd_sc_hd__inv_2 \inv[67]/_0_  (.A(\inv_in[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[68] ));
 sky130_fd_sc_hd__inv_2 \inv[680]/_0_  (.A(\inv_in[680] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[681] ));
 sky130_fd_sc_hd__inv_2 \inv[681]/_0_  (.A(\inv_in[681] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[682] ));
 sky130_fd_sc_hd__inv_2 \inv[682]/_0_  (.A(\inv_in[682] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[683] ));
 sky130_fd_sc_hd__inv_2 \inv[683]/_0_  (.A(\inv_in[683] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[684] ));
 sky130_fd_sc_hd__inv_2 \inv[684]/_0_  (.A(\inv_in[684] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[685] ));
 sky130_fd_sc_hd__inv_2 \inv[685]/_0_  (.A(\inv_in[685] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[686] ));
 sky130_fd_sc_hd__inv_2 \inv[686]/_0_  (.A(\inv_in[686] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[687] ));
 sky130_fd_sc_hd__inv_2 \inv[687]/_0_  (.A(\inv_in[687] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[688] ));
 sky130_fd_sc_hd__inv_2 \inv[688]/_0_  (.A(\inv_in[688] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[689] ));
 sky130_fd_sc_hd__inv_2 \inv[689]/_0_  (.A(\inv_in[689] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[690] ));
 sky130_fd_sc_hd__inv_2 \inv[68]/_0_  (.A(\inv_in[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[69] ));
 sky130_fd_sc_hd__inv_2 \inv[690]/_0_  (.A(\inv_in[690] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[691] ));
 sky130_fd_sc_hd__inv_2 \inv[691]/_0_  (.A(\inv_in[691] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[692] ));
 sky130_fd_sc_hd__inv_2 \inv[692]/_0_  (.A(\inv_in[692] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[693] ));
 sky130_fd_sc_hd__inv_2 \inv[693]/_0_  (.A(\inv_in[693] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[694] ));
 sky130_fd_sc_hd__inv_2 \inv[694]/_0_  (.A(\inv_in[694] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[695] ));
 sky130_fd_sc_hd__inv_2 \inv[695]/_0_  (.A(\inv_in[695] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[696] ));
 sky130_fd_sc_hd__inv_2 \inv[696]/_0_  (.A(\inv_in[696] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[697] ));
 sky130_fd_sc_hd__inv_2 \inv[697]/_0_  (.A(\inv_in[697] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[698] ));
 sky130_fd_sc_hd__inv_2 \inv[698]/_0_  (.A(\inv_in[698] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[699] ));
 sky130_fd_sc_hd__inv_2 \inv[699]/_0_  (.A(\inv_in[699] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[700] ));
 sky130_fd_sc_hd__inv_2 \inv[69]/_0_  (.A(\inv_in[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[70] ));
 sky130_fd_sc_hd__inv_2 \inv[6]/_0_  (.A(\inv_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[7] ));
 sky130_fd_sc_hd__inv_2 \inv[700]/_0_  (.A(\inv_in[700] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[701] ));
 sky130_fd_sc_hd__inv_2 \inv[701]/_0_  (.A(\inv_in[701] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[702] ));
 sky130_fd_sc_hd__inv_2 \inv[702]/_0_  (.A(\inv_in[702] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[703] ));
 sky130_fd_sc_hd__inv_2 \inv[703]/_0_  (.A(\inv_in[703] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[704] ));
 sky130_fd_sc_hd__inv_2 \inv[704]/_0_  (.A(\inv_in[704] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[705] ));
 sky130_fd_sc_hd__inv_2 \inv[705]/_0_  (.A(\inv_in[705] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[706] ));
 sky130_fd_sc_hd__inv_2 \inv[706]/_0_  (.A(\inv_in[706] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[707] ));
 sky130_fd_sc_hd__inv_2 \inv[707]/_0_  (.A(\inv_in[707] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[708] ));
 sky130_fd_sc_hd__inv_2 \inv[708]/_0_  (.A(\inv_in[708] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[709] ));
 sky130_fd_sc_hd__inv_2 \inv[709]/_0_  (.A(\inv_in[709] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[710] ));
 sky130_fd_sc_hd__inv_2 \inv[70]/_0_  (.A(\inv_in[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[71] ));
 sky130_fd_sc_hd__inv_2 \inv[710]/_0_  (.A(\inv_in[710] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[711] ));
 sky130_fd_sc_hd__inv_2 \inv[711]/_0_  (.A(\inv_in[711] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[712] ));
 sky130_fd_sc_hd__inv_2 \inv[712]/_0_  (.A(\inv_in[712] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[713] ));
 sky130_fd_sc_hd__inv_2 \inv[713]/_0_  (.A(\inv_in[713] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[714] ));
 sky130_fd_sc_hd__inv_2 \inv[714]/_0_  (.A(\inv_in[714] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[715] ));
 sky130_fd_sc_hd__inv_2 \inv[715]/_0_  (.A(\inv_in[715] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[716] ));
 sky130_fd_sc_hd__inv_2 \inv[716]/_0_  (.A(\inv_in[716] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[717] ));
 sky130_fd_sc_hd__inv_2 \inv[717]/_0_  (.A(\inv_in[717] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[718] ));
 sky130_fd_sc_hd__inv_2 \inv[718]/_0_  (.A(\inv_in[718] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[719] ));
 sky130_fd_sc_hd__inv_2 \inv[719]/_0_  (.A(\inv_in[719] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[720] ));
 sky130_fd_sc_hd__inv_2 \inv[71]/_0_  (.A(\inv_in[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[72] ));
 sky130_fd_sc_hd__inv_2 \inv[720]/_0_  (.A(\inv_in[720] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[721] ));
 sky130_fd_sc_hd__inv_2 \inv[721]/_0_  (.A(\inv_in[721] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[722] ));
 sky130_fd_sc_hd__inv_2 \inv[722]/_0_  (.A(\inv_in[722] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[723] ));
 sky130_fd_sc_hd__inv_2 \inv[723]/_0_  (.A(\inv_in[723] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[724] ));
 sky130_fd_sc_hd__inv_2 \inv[724]/_0_  (.A(\inv_in[724] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[725] ));
 sky130_fd_sc_hd__inv_2 \inv[725]/_0_  (.A(\inv_in[725] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[726] ));
 sky130_fd_sc_hd__inv_2 \inv[726]/_0_  (.A(\inv_in[726] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[727] ));
 sky130_fd_sc_hd__inv_2 \inv[727]/_0_  (.A(\inv_in[727] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[728] ));
 sky130_fd_sc_hd__inv_2 \inv[728]/_0_  (.A(\inv_in[728] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[729] ));
 sky130_fd_sc_hd__inv_2 \inv[729]/_0_  (.A(\inv_in[729] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[730] ));
 sky130_fd_sc_hd__inv_2 \inv[72]/_0_  (.A(\inv_in[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[73] ));
 sky130_fd_sc_hd__inv_2 \inv[730]/_0_  (.A(\inv_in[730] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[731] ));
 sky130_fd_sc_hd__inv_2 \inv[731]/_0_  (.A(\inv_in[731] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[732] ));
 sky130_fd_sc_hd__inv_2 \inv[732]/_0_  (.A(\inv_in[732] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[733] ));
 sky130_fd_sc_hd__inv_2 \inv[733]/_0_  (.A(\inv_in[733] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[734] ));
 sky130_fd_sc_hd__inv_2 \inv[734]/_0_  (.A(\inv_in[734] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[735] ));
 sky130_fd_sc_hd__inv_2 \inv[735]/_0_  (.A(\inv_in[735] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[736] ));
 sky130_fd_sc_hd__inv_2 \inv[736]/_0_  (.A(\inv_in[736] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[737] ));
 sky130_fd_sc_hd__inv_2 \inv[737]/_0_  (.A(\inv_in[737] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[738] ));
 sky130_fd_sc_hd__inv_2 \inv[738]/_0_  (.A(\inv_in[738] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[739] ));
 sky130_fd_sc_hd__inv_2 \inv[739]/_0_  (.A(\inv_in[739] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[740] ));
 sky130_fd_sc_hd__inv_2 \inv[73]/_0_  (.A(\inv_in[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[74] ));
 sky130_fd_sc_hd__inv_2 \inv[740]/_0_  (.A(\inv_in[740] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[741] ));
 sky130_fd_sc_hd__inv_2 \inv[741]/_0_  (.A(\inv_in[741] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[742] ));
 sky130_fd_sc_hd__inv_2 \inv[742]/_0_  (.A(\inv_in[742] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[743] ));
 sky130_fd_sc_hd__inv_2 \inv[743]/_0_  (.A(\inv_in[743] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[744] ));
 sky130_fd_sc_hd__inv_2 \inv[744]/_0_  (.A(\inv_in[744] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[745] ));
 sky130_fd_sc_hd__inv_2 \inv[745]/_0_  (.A(\inv_in[745] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[746] ));
 sky130_fd_sc_hd__inv_2 \inv[746]/_0_  (.A(\inv_in[746] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[747] ));
 sky130_fd_sc_hd__inv_2 \inv[747]/_0_  (.A(\inv_in[747] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[748] ));
 sky130_fd_sc_hd__inv_2 \inv[748]/_0_  (.A(\inv_in[748] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[749] ));
 sky130_fd_sc_hd__inv_2 \inv[749]/_0_  (.A(\inv_in[749] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[750] ));
 sky130_fd_sc_hd__inv_2 \inv[74]/_0_  (.A(\inv_in[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[75] ));
 sky130_fd_sc_hd__inv_2 \inv[750]/_0_  (.A(\inv_in[750] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[751] ));
 sky130_fd_sc_hd__inv_2 \inv[751]/_0_  (.A(\inv_in[751] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[752] ));
 sky130_fd_sc_hd__inv_2 \inv[752]/_0_  (.A(\inv_in[752] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[753] ));
 sky130_fd_sc_hd__inv_2 \inv[753]/_0_  (.A(\inv_in[753] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[754] ));
 sky130_fd_sc_hd__inv_2 \inv[754]/_0_  (.A(\inv_in[754] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[755] ));
 sky130_fd_sc_hd__inv_2 \inv[755]/_0_  (.A(\inv_in[755] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[756] ));
 sky130_fd_sc_hd__inv_2 \inv[756]/_0_  (.A(\inv_in[756] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[757] ));
 sky130_fd_sc_hd__inv_2 \inv[757]/_0_  (.A(\inv_in[757] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[758] ));
 sky130_fd_sc_hd__inv_2 \inv[758]/_0_  (.A(\inv_in[758] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[759] ));
 sky130_fd_sc_hd__inv_2 \inv[759]/_0_  (.A(\inv_in[759] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[760] ));
 sky130_fd_sc_hd__inv_2 \inv[75]/_0_  (.A(\inv_in[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[76] ));
 sky130_fd_sc_hd__inv_2 \inv[760]/_0_  (.A(\inv_in[760] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[761] ));
 sky130_fd_sc_hd__inv_2 \inv[761]/_0_  (.A(\inv_in[761] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[762] ));
 sky130_fd_sc_hd__inv_2 \inv[762]/_0_  (.A(\inv_in[762] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[763] ));
 sky130_fd_sc_hd__inv_2 \inv[763]/_0_  (.A(\inv_in[763] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[764] ));
 sky130_fd_sc_hd__inv_2 \inv[764]/_0_  (.A(\inv_in[764] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[765] ));
 sky130_fd_sc_hd__inv_2 \inv[765]/_0_  (.A(\inv_in[765] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[766] ));
 sky130_fd_sc_hd__inv_2 \inv[766]/_0_  (.A(\inv_in[766] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[767] ));
 sky130_fd_sc_hd__inv_2 \inv[767]/_0_  (.A(\inv_in[767] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[768] ));
 sky130_fd_sc_hd__inv_2 \inv[768]/_0_  (.A(\inv_in[768] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[769] ));
 sky130_fd_sc_hd__inv_2 \inv[769]/_0_  (.A(\inv_in[769] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[770] ));
 sky130_fd_sc_hd__inv_2 \inv[76]/_0_  (.A(\inv_in[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[77] ));
 sky130_fd_sc_hd__inv_2 \inv[770]/_0_  (.A(\inv_in[770] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[771] ));
 sky130_fd_sc_hd__inv_2 \inv[771]/_0_  (.A(\inv_in[771] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[772] ));
 sky130_fd_sc_hd__inv_2 \inv[772]/_0_  (.A(\inv_in[772] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[773] ));
 sky130_fd_sc_hd__inv_2 \inv[773]/_0_  (.A(\inv_in[773] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[774] ));
 sky130_fd_sc_hd__inv_2 \inv[774]/_0_  (.A(\inv_in[774] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[775] ));
 sky130_fd_sc_hd__inv_2 \inv[775]/_0_  (.A(\inv_in[775] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[776] ));
 sky130_fd_sc_hd__inv_2 \inv[776]/_0_  (.A(\inv_in[776] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[777] ));
 sky130_fd_sc_hd__inv_2 \inv[777]/_0_  (.A(\inv_in[777] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[778] ));
 sky130_fd_sc_hd__inv_2 \inv[778]/_0_  (.A(\inv_in[778] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[779] ));
 sky130_fd_sc_hd__inv_2 \inv[779]/_0_  (.A(\inv_in[779] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[780] ));
 sky130_fd_sc_hd__inv_2 \inv[77]/_0_  (.A(\inv_in[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[78] ));
 sky130_fd_sc_hd__inv_2 \inv[780]/_0_  (.A(\inv_in[780] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[781] ));
 sky130_fd_sc_hd__inv_2 \inv[781]/_0_  (.A(\inv_in[781] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[782] ));
 sky130_fd_sc_hd__inv_2 \inv[782]/_0_  (.A(\inv_in[782] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[783] ));
 sky130_fd_sc_hd__inv_2 \inv[783]/_0_  (.A(\inv_in[783] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[784] ));
 sky130_fd_sc_hd__inv_2 \inv[784]/_0_  (.A(\inv_in[784] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[785] ));
 sky130_fd_sc_hd__inv_2 \inv[785]/_0_  (.A(\inv_in[785] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[786] ));
 sky130_fd_sc_hd__inv_2 \inv[786]/_0_  (.A(\inv_in[786] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[787] ));
 sky130_fd_sc_hd__inv_2 \inv[787]/_0_  (.A(\inv_in[787] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[788] ));
 sky130_fd_sc_hd__inv_2 \inv[788]/_0_  (.A(\inv_in[788] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[789] ));
 sky130_fd_sc_hd__inv_2 \inv[789]/_0_  (.A(\inv_in[789] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[790] ));
 sky130_fd_sc_hd__inv_2 \inv[78]/_0_  (.A(\inv_in[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[79] ));
 sky130_fd_sc_hd__inv_2 \inv[790]/_0_  (.A(\inv_in[790] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[791] ));
 sky130_fd_sc_hd__inv_2 \inv[791]/_0_  (.A(\inv_in[791] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[792] ));
 sky130_fd_sc_hd__inv_2 \inv[792]/_0_  (.A(\inv_in[792] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[793] ));
 sky130_fd_sc_hd__inv_2 \inv[793]/_0_  (.A(\inv_in[793] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[794] ));
 sky130_fd_sc_hd__inv_2 \inv[794]/_0_  (.A(\inv_in[794] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[795] ));
 sky130_fd_sc_hd__inv_2 \inv[795]/_0_  (.A(\inv_in[795] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[796] ));
 sky130_fd_sc_hd__inv_2 \inv[796]/_0_  (.A(\inv_in[796] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[797] ));
 sky130_fd_sc_hd__inv_2 \inv[797]/_0_  (.A(\inv_in[797] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[798] ));
 sky130_fd_sc_hd__inv_2 \inv[798]/_0_  (.A(\inv_in[798] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[799] ));
 sky130_fd_sc_hd__inv_2 \inv[799]/_0_  (.A(\inv_in[799] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[800] ));
 sky130_fd_sc_hd__inv_2 \inv[79]/_0_  (.A(\inv_in[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[80] ));
 sky130_fd_sc_hd__inv_2 \inv[7]/_0_  (.A(\inv_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[8] ));
 sky130_fd_sc_hd__inv_2 \inv[800]/_0_  (.A(\inv_in[800] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[801] ));
 sky130_fd_sc_hd__inv_2 \inv[801]/_0_  (.A(\inv_in[801] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[802] ));
 sky130_fd_sc_hd__inv_2 \inv[802]/_0_  (.A(\inv_in[802] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[803] ));
 sky130_fd_sc_hd__inv_2 \inv[803]/_0_  (.A(\inv_in[803] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[804] ));
 sky130_fd_sc_hd__inv_2 \inv[804]/_0_  (.A(\inv_in[804] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[805] ));
 sky130_fd_sc_hd__inv_2 \inv[805]/_0_  (.A(\inv_in[805] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[806] ));
 sky130_fd_sc_hd__inv_2 \inv[806]/_0_  (.A(\inv_in[806] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[807] ));
 sky130_fd_sc_hd__inv_2 \inv[807]/_0_  (.A(\inv_in[807] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[808] ));
 sky130_fd_sc_hd__inv_2 \inv[808]/_0_  (.A(\inv_in[808] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[809] ));
 sky130_fd_sc_hd__inv_2 \inv[809]/_0_  (.A(\inv_in[809] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[810] ));
 sky130_fd_sc_hd__inv_2 \inv[80]/_0_  (.A(\inv_in[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[81] ));
 sky130_fd_sc_hd__inv_2 \inv[810]/_0_  (.A(\inv_in[810] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[811] ));
 sky130_fd_sc_hd__inv_2 \inv[811]/_0_  (.A(\inv_in[811] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[812] ));
 sky130_fd_sc_hd__inv_2 \inv[812]/_0_  (.A(\inv_in[812] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[813] ));
 sky130_fd_sc_hd__inv_2 \inv[813]/_0_  (.A(\inv_in[813] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[814] ));
 sky130_fd_sc_hd__inv_2 \inv[814]/_0_  (.A(\inv_in[814] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[815] ));
 sky130_fd_sc_hd__inv_2 \inv[815]/_0_  (.A(\inv_in[815] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[816] ));
 sky130_fd_sc_hd__inv_2 \inv[816]/_0_  (.A(\inv_in[816] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[817] ));
 sky130_fd_sc_hd__inv_2 \inv[817]/_0_  (.A(\inv_in[817] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[818] ));
 sky130_fd_sc_hd__inv_2 \inv[818]/_0_  (.A(\inv_in[818] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[819] ));
 sky130_fd_sc_hd__inv_2 \inv[819]/_0_  (.A(\inv_in[819] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[820] ));
 sky130_fd_sc_hd__inv_2 \inv[81]/_0_  (.A(\inv_in[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[82] ));
 sky130_fd_sc_hd__inv_2 \inv[820]/_0_  (.A(\inv_in[820] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[821] ));
 sky130_fd_sc_hd__inv_2 \inv[821]/_0_  (.A(\inv_in[821] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[822] ));
 sky130_fd_sc_hd__inv_2 \inv[822]/_0_  (.A(\inv_in[822] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[823] ));
 sky130_fd_sc_hd__inv_2 \inv[823]/_0_  (.A(\inv_in[823] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[824] ));
 sky130_fd_sc_hd__inv_2 \inv[824]/_0_  (.A(\inv_in[824] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[825] ));
 sky130_fd_sc_hd__inv_2 \inv[825]/_0_  (.A(\inv_in[825] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[826] ));
 sky130_fd_sc_hd__inv_2 \inv[826]/_0_  (.A(\inv_in[826] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[827] ));
 sky130_fd_sc_hd__inv_2 \inv[827]/_0_  (.A(\inv_in[827] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[828] ));
 sky130_fd_sc_hd__inv_2 \inv[828]/_0_  (.A(\inv_in[828] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[829] ));
 sky130_fd_sc_hd__inv_2 \inv[829]/_0_  (.A(\inv_in[829] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[830] ));
 sky130_fd_sc_hd__inv_2 \inv[82]/_0_  (.A(\inv_in[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[83] ));
 sky130_fd_sc_hd__inv_2 \inv[830]/_0_  (.A(\inv_in[830] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[831] ));
 sky130_fd_sc_hd__inv_2 \inv[831]/_0_  (.A(\inv_in[831] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[832] ));
 sky130_fd_sc_hd__inv_2 \inv[832]/_0_  (.A(\inv_in[832] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[833] ));
 sky130_fd_sc_hd__inv_2 \inv[833]/_0_  (.A(\inv_in[833] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[834] ));
 sky130_fd_sc_hd__inv_2 \inv[834]/_0_  (.A(\inv_in[834] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[835] ));
 sky130_fd_sc_hd__inv_2 \inv[835]/_0_  (.A(\inv_in[835] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[836] ));
 sky130_fd_sc_hd__inv_2 \inv[836]/_0_  (.A(\inv_in[836] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[837] ));
 sky130_fd_sc_hd__inv_2 \inv[837]/_0_  (.A(\inv_in[837] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[838] ));
 sky130_fd_sc_hd__inv_2 \inv[838]/_0_  (.A(\inv_in[838] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[839] ));
 sky130_fd_sc_hd__inv_2 \inv[839]/_0_  (.A(\inv_in[839] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[840] ));
 sky130_fd_sc_hd__inv_2 \inv[83]/_0_  (.A(\inv_in[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[84] ));
 sky130_fd_sc_hd__inv_2 \inv[840]/_0_  (.A(\inv_in[840] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[841] ));
 sky130_fd_sc_hd__inv_2 \inv[841]/_0_  (.A(\inv_in[841] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[842] ));
 sky130_fd_sc_hd__inv_2 \inv[842]/_0_  (.A(\inv_in[842] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[843] ));
 sky130_fd_sc_hd__inv_2 \inv[843]/_0_  (.A(\inv_in[843] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[844] ));
 sky130_fd_sc_hd__inv_2 \inv[844]/_0_  (.A(\inv_in[844] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[845] ));
 sky130_fd_sc_hd__inv_2 \inv[845]/_0_  (.A(\inv_in[845] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[846] ));
 sky130_fd_sc_hd__inv_2 \inv[846]/_0_  (.A(\inv_in[846] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[847] ));
 sky130_fd_sc_hd__inv_2 \inv[847]/_0_  (.A(\inv_in[847] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[848] ));
 sky130_fd_sc_hd__inv_2 \inv[848]/_0_  (.A(\inv_in[848] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[849] ));
 sky130_fd_sc_hd__inv_2 \inv[849]/_0_  (.A(\inv_in[849] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[850] ));
 sky130_fd_sc_hd__inv_2 \inv[84]/_0_  (.A(\inv_in[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[85] ));
 sky130_fd_sc_hd__inv_2 \inv[850]/_0_  (.A(\inv_in[850] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[851] ));
 sky130_fd_sc_hd__inv_2 \inv[851]/_0_  (.A(\inv_in[851] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[852] ));
 sky130_fd_sc_hd__inv_2 \inv[852]/_0_  (.A(\inv_in[852] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[853] ));
 sky130_fd_sc_hd__inv_2 \inv[853]/_0_  (.A(\inv_in[853] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[854] ));
 sky130_fd_sc_hd__inv_2 \inv[854]/_0_  (.A(\inv_in[854] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[855] ));
 sky130_fd_sc_hd__inv_2 \inv[855]/_0_  (.A(\inv_in[855] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[856] ));
 sky130_fd_sc_hd__inv_2 \inv[856]/_0_  (.A(\inv_in[856] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[857] ));
 sky130_fd_sc_hd__inv_2 \inv[857]/_0_  (.A(\inv_in[857] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[858] ));
 sky130_fd_sc_hd__inv_2 \inv[858]/_0_  (.A(\inv_in[858] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[859] ));
 sky130_fd_sc_hd__inv_2 \inv[859]/_0_  (.A(\inv_in[859] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[860] ));
 sky130_fd_sc_hd__inv_2 \inv[85]/_0_  (.A(\inv_in[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[86] ));
 sky130_fd_sc_hd__inv_2 \inv[860]/_0_  (.A(\inv_in[860] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[861] ));
 sky130_fd_sc_hd__inv_2 \inv[861]/_0_  (.A(\inv_in[861] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[862] ));
 sky130_fd_sc_hd__inv_2 \inv[862]/_0_  (.A(\inv_in[862] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[863] ));
 sky130_fd_sc_hd__inv_2 \inv[863]/_0_  (.A(\inv_in[863] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[864] ));
 sky130_fd_sc_hd__inv_2 \inv[864]/_0_  (.A(\inv_in[864] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[865] ));
 sky130_fd_sc_hd__inv_2 \inv[865]/_0_  (.A(\inv_in[865] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[866] ));
 sky130_fd_sc_hd__inv_2 \inv[866]/_0_  (.A(\inv_in[866] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[867] ));
 sky130_fd_sc_hd__inv_2 \inv[867]/_0_  (.A(\inv_in[867] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[868] ));
 sky130_fd_sc_hd__inv_2 \inv[868]/_0_  (.A(\inv_in[868] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[869] ));
 sky130_fd_sc_hd__inv_2 \inv[869]/_0_  (.A(\inv_in[869] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[870] ));
 sky130_fd_sc_hd__inv_2 \inv[86]/_0_  (.A(\inv_in[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[87] ));
 sky130_fd_sc_hd__inv_2 \inv[870]/_0_  (.A(\inv_in[870] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[871] ));
 sky130_fd_sc_hd__inv_2 \inv[871]/_0_  (.A(\inv_in[871] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[872] ));
 sky130_fd_sc_hd__inv_2 \inv[872]/_0_  (.A(\inv_in[872] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[873] ));
 sky130_fd_sc_hd__inv_2 \inv[873]/_0_  (.A(\inv_in[873] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[874] ));
 sky130_fd_sc_hd__inv_2 \inv[874]/_0_  (.A(\inv_in[874] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[875] ));
 sky130_fd_sc_hd__inv_2 \inv[875]/_0_  (.A(\inv_in[875] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[876] ));
 sky130_fd_sc_hd__inv_2 \inv[876]/_0_  (.A(\inv_in[876] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[877] ));
 sky130_fd_sc_hd__inv_2 \inv[877]/_0_  (.A(\inv_in[877] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[878] ));
 sky130_fd_sc_hd__inv_2 \inv[878]/_0_  (.A(\inv_in[878] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[879] ));
 sky130_fd_sc_hd__inv_2 \inv[879]/_0_  (.A(\inv_in[879] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[880] ));
 sky130_fd_sc_hd__inv_2 \inv[87]/_0_  (.A(\inv_in[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[88] ));
 sky130_fd_sc_hd__inv_2 \inv[880]/_0_  (.A(\inv_in[880] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[881] ));
 sky130_fd_sc_hd__inv_2 \inv[881]/_0_  (.A(\inv_in[881] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[882] ));
 sky130_fd_sc_hd__inv_2 \inv[882]/_0_  (.A(\inv_in[882] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[883] ));
 sky130_fd_sc_hd__inv_2 \inv[883]/_0_  (.A(\inv_in[883] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[884] ));
 sky130_fd_sc_hd__inv_2 \inv[884]/_0_  (.A(\inv_in[884] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[885] ));
 sky130_fd_sc_hd__inv_2 \inv[885]/_0_  (.A(\inv_in[885] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[886] ));
 sky130_fd_sc_hd__inv_2 \inv[886]/_0_  (.A(\inv_in[886] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[887] ));
 sky130_fd_sc_hd__inv_2 \inv[887]/_0_  (.A(\inv_in[887] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[888] ));
 sky130_fd_sc_hd__inv_2 \inv[888]/_0_  (.A(\inv_in[888] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[889] ));
 sky130_fd_sc_hd__inv_2 \inv[889]/_0_  (.A(\inv_in[889] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[890] ));
 sky130_fd_sc_hd__inv_2 \inv[88]/_0_  (.A(\inv_in[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[89] ));
 sky130_fd_sc_hd__inv_2 \inv[890]/_0_  (.A(\inv_in[890] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[891] ));
 sky130_fd_sc_hd__inv_2 \inv[891]/_0_  (.A(\inv_in[891] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[892] ));
 sky130_fd_sc_hd__inv_2 \inv[892]/_0_  (.A(\inv_in[892] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[893] ));
 sky130_fd_sc_hd__inv_2 \inv[893]/_0_  (.A(\inv_in[893] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[894] ));
 sky130_fd_sc_hd__inv_2 \inv[894]/_0_  (.A(\inv_in[894] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[895] ));
 sky130_fd_sc_hd__inv_2 \inv[895]/_0_  (.A(\inv_in[895] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[896] ));
 sky130_fd_sc_hd__inv_2 \inv[896]/_0_  (.A(\inv_in[896] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[897] ));
 sky130_fd_sc_hd__inv_2 \inv[897]/_0_  (.A(\inv_in[897] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[898] ));
 sky130_fd_sc_hd__inv_2 \inv[898]/_0_  (.A(\inv_in[898] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[899] ));
 sky130_fd_sc_hd__inv_2 \inv[899]/_0_  (.A(\inv_in[899] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[900] ));
 sky130_fd_sc_hd__inv_2 \inv[89]/_0_  (.A(\inv_in[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[90] ));
 sky130_fd_sc_hd__inv_2 \inv[8]/_0_  (.A(\inv_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[9] ));
 sky130_fd_sc_hd__inv_2 \inv[900]/_0_  (.A(\inv_in[900] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[901] ));
 sky130_fd_sc_hd__inv_2 \inv[901]/_0_  (.A(\inv_in[901] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[902] ));
 sky130_fd_sc_hd__inv_2 \inv[902]/_0_  (.A(\inv_in[902] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[903] ));
 sky130_fd_sc_hd__inv_2 \inv[903]/_0_  (.A(\inv_in[903] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[904] ));
 sky130_fd_sc_hd__inv_2 \inv[904]/_0_  (.A(\inv_in[904] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[905] ));
 sky130_fd_sc_hd__inv_2 \inv[905]/_0_  (.A(\inv_in[905] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[906] ));
 sky130_fd_sc_hd__inv_2 \inv[906]/_0_  (.A(\inv_in[906] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[907] ));
 sky130_fd_sc_hd__inv_2 \inv[907]/_0_  (.A(\inv_in[907] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[908] ));
 sky130_fd_sc_hd__inv_2 \inv[908]/_0_  (.A(\inv_in[908] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[909] ));
 sky130_fd_sc_hd__inv_2 \inv[909]/_0_  (.A(\inv_in[909] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[910] ));
 sky130_fd_sc_hd__inv_2 \inv[90]/_0_  (.A(\inv_in[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[91] ));
 sky130_fd_sc_hd__inv_2 \inv[910]/_0_  (.A(\inv_in[910] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[911] ));
 sky130_fd_sc_hd__inv_2 \inv[911]/_0_  (.A(\inv_in[911] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[912] ));
 sky130_fd_sc_hd__inv_2 \inv[912]/_0_  (.A(\inv_in[912] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[913] ));
 sky130_fd_sc_hd__inv_2 \inv[913]/_0_  (.A(\inv_in[913] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[914] ));
 sky130_fd_sc_hd__inv_2 \inv[914]/_0_  (.A(\inv_in[914] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[915] ));
 sky130_fd_sc_hd__inv_2 \inv[915]/_0_  (.A(\inv_in[915] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[916] ));
 sky130_fd_sc_hd__inv_2 \inv[916]/_0_  (.A(\inv_in[916] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[917] ));
 sky130_fd_sc_hd__inv_2 \inv[917]/_0_  (.A(\inv_in[917] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[918] ));
 sky130_fd_sc_hd__inv_2 \inv[918]/_0_  (.A(\inv_in[918] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[919] ));
 sky130_fd_sc_hd__inv_2 \inv[919]/_0_  (.A(\inv_in[919] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[920] ));
 sky130_fd_sc_hd__inv_2 \inv[91]/_0_  (.A(\inv_in[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[92] ));
 sky130_fd_sc_hd__inv_2 \inv[920]/_0_  (.A(\inv_in[920] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[921] ));
 sky130_fd_sc_hd__inv_2 \inv[921]/_0_  (.A(\inv_in[921] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[922] ));
 sky130_fd_sc_hd__inv_2 \inv[922]/_0_  (.A(\inv_in[922] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[923] ));
 sky130_fd_sc_hd__inv_2 \inv[923]/_0_  (.A(\inv_in[923] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[924] ));
 sky130_fd_sc_hd__inv_2 \inv[924]/_0_  (.A(\inv_in[924] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[925] ));
 sky130_fd_sc_hd__inv_2 \inv[925]/_0_  (.A(\inv_in[925] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[926] ));
 sky130_fd_sc_hd__inv_2 \inv[926]/_0_  (.A(\inv_in[926] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[927] ));
 sky130_fd_sc_hd__inv_2 \inv[927]/_0_  (.A(\inv_in[927] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[928] ));
 sky130_fd_sc_hd__inv_2 \inv[928]/_0_  (.A(\inv_in[928] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[929] ));
 sky130_fd_sc_hd__inv_2 \inv[929]/_0_  (.A(\inv_in[929] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[930] ));
 sky130_fd_sc_hd__inv_2 \inv[92]/_0_  (.A(\inv_in[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[93] ));
 sky130_fd_sc_hd__inv_2 \inv[930]/_0_  (.A(\inv_in[930] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[931] ));
 sky130_fd_sc_hd__inv_2 \inv[931]/_0_  (.A(\inv_in[931] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[932] ));
 sky130_fd_sc_hd__inv_2 \inv[932]/_0_  (.A(\inv_in[932] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[933] ));
 sky130_fd_sc_hd__inv_2 \inv[933]/_0_  (.A(\inv_in[933] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[934] ));
 sky130_fd_sc_hd__inv_2 \inv[934]/_0_  (.A(\inv_in[934] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[935] ));
 sky130_fd_sc_hd__inv_2 \inv[935]/_0_  (.A(\inv_in[935] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[936] ));
 sky130_fd_sc_hd__inv_2 \inv[936]/_0_  (.A(\inv_in[936] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[937] ));
 sky130_fd_sc_hd__inv_2 \inv[937]/_0_  (.A(\inv_in[937] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[938] ));
 sky130_fd_sc_hd__inv_2 \inv[938]/_0_  (.A(\inv_in[938] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[939] ));
 sky130_fd_sc_hd__inv_2 \inv[939]/_0_  (.A(\inv_in[939] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[940] ));
 sky130_fd_sc_hd__inv_2 \inv[93]/_0_  (.A(\inv_in[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[94] ));
 sky130_fd_sc_hd__inv_2 \inv[940]/_0_  (.A(\inv_in[940] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[941] ));
 sky130_fd_sc_hd__inv_2 \inv[941]/_0_  (.A(\inv_in[941] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[942] ));
 sky130_fd_sc_hd__inv_2 \inv[942]/_0_  (.A(\inv_in[942] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[943] ));
 sky130_fd_sc_hd__inv_2 \inv[943]/_0_  (.A(\inv_in[943] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[944] ));
 sky130_fd_sc_hd__inv_2 \inv[944]/_0_  (.A(\inv_in[944] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[945] ));
 sky130_fd_sc_hd__inv_2 \inv[945]/_0_  (.A(\inv_in[945] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[946] ));
 sky130_fd_sc_hd__inv_2 \inv[946]/_0_  (.A(\inv_in[946] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[947] ));
 sky130_fd_sc_hd__inv_2 \inv[947]/_0_  (.A(\inv_in[947] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[948] ));
 sky130_fd_sc_hd__inv_2 \inv[948]/_0_  (.A(\inv_in[948] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[949] ));
 sky130_fd_sc_hd__inv_2 \inv[949]/_0_  (.A(\inv_in[949] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[950] ));
 sky130_fd_sc_hd__inv_2 \inv[94]/_0_  (.A(\inv_in[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[95] ));
 sky130_fd_sc_hd__inv_2 \inv[950]/_0_  (.A(\inv_in[950] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[951] ));
 sky130_fd_sc_hd__inv_2 \inv[951]/_0_  (.A(\inv_in[951] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[952] ));
 sky130_fd_sc_hd__inv_2 \inv[952]/_0_  (.A(\inv_in[952] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[953] ));
 sky130_fd_sc_hd__inv_2 \inv[953]/_0_  (.A(\inv_in[953] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[954] ));
 sky130_fd_sc_hd__inv_2 \inv[954]/_0_  (.A(\inv_in[954] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[955] ));
 sky130_fd_sc_hd__inv_2 \inv[955]/_0_  (.A(\inv_in[955] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[956] ));
 sky130_fd_sc_hd__inv_2 \inv[956]/_0_  (.A(\inv_in[956] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[957] ));
 sky130_fd_sc_hd__inv_2 \inv[957]/_0_  (.A(\inv_in[957] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[958] ));
 sky130_fd_sc_hd__inv_2 \inv[958]/_0_  (.A(\inv_in[958] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[959] ));
 sky130_fd_sc_hd__inv_2 \inv[959]/_0_  (.A(\inv_in[959] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[960] ));
 sky130_fd_sc_hd__inv_2 \inv[95]/_0_  (.A(\inv_in[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[96] ));
 sky130_fd_sc_hd__inv_2 \inv[960]/_0_  (.A(\inv_in[960] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[961] ));
 sky130_fd_sc_hd__inv_2 \inv[961]/_0_  (.A(\inv_in[961] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[962] ));
 sky130_fd_sc_hd__inv_2 \inv[962]/_0_  (.A(\inv_in[962] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[963] ));
 sky130_fd_sc_hd__inv_2 \inv[963]/_0_  (.A(\inv_in[963] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[964] ));
 sky130_fd_sc_hd__inv_2 \inv[964]/_0_  (.A(\inv_in[964] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[965] ));
 sky130_fd_sc_hd__inv_2 \inv[965]/_0_  (.A(\inv_in[965] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[966] ));
 sky130_fd_sc_hd__inv_2 \inv[966]/_0_  (.A(\inv_in[966] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[967] ));
 sky130_fd_sc_hd__inv_2 \inv[967]/_0_  (.A(\inv_in[967] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[968] ));
 sky130_fd_sc_hd__inv_2 \inv[968]/_0_  (.A(\inv_in[968] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[969] ));
 sky130_fd_sc_hd__inv_2 \inv[969]/_0_  (.A(\inv_in[969] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[970] ));
 sky130_fd_sc_hd__inv_2 \inv[96]/_0_  (.A(\inv_in[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[97] ));
 sky130_fd_sc_hd__inv_2 \inv[970]/_0_  (.A(\inv_in[970] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[971] ));
 sky130_fd_sc_hd__inv_2 \inv[971]/_0_  (.A(\inv_in[971] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[972] ));
 sky130_fd_sc_hd__inv_2 \inv[972]/_0_  (.A(\inv_in[972] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[973] ));
 sky130_fd_sc_hd__inv_2 \inv[973]/_0_  (.A(\inv_in[973] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[974] ));
 sky130_fd_sc_hd__inv_2 \inv[974]/_0_  (.A(\inv_in[974] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[975] ));
 sky130_fd_sc_hd__inv_2 \inv[975]/_0_  (.A(\inv_in[975] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[976] ));
 sky130_fd_sc_hd__inv_2 \inv[976]/_0_  (.A(\inv_in[976] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[977] ));
 sky130_fd_sc_hd__inv_2 \inv[977]/_0_  (.A(\inv_in[977] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[978] ));
 sky130_fd_sc_hd__inv_2 \inv[978]/_0_  (.A(\inv_in[978] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[979] ));
 sky130_fd_sc_hd__inv_2 \inv[979]/_0_  (.A(\inv_in[979] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[980] ));
 sky130_fd_sc_hd__inv_2 \inv[97]/_0_  (.A(\inv_in[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[98] ));
 sky130_fd_sc_hd__inv_2 \inv[980]/_0_  (.A(\inv_in[980] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[981] ));
 sky130_fd_sc_hd__inv_2 \inv[981]/_0_  (.A(\inv_in[981] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[982] ));
 sky130_fd_sc_hd__inv_2 \inv[982]/_0_  (.A(\inv_in[982] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[983] ));
 sky130_fd_sc_hd__inv_2 \inv[983]/_0_  (.A(\inv_in[983] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[984] ));
 sky130_fd_sc_hd__inv_2 \inv[984]/_0_  (.A(\inv_in[984] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[985] ));
 sky130_fd_sc_hd__inv_2 \inv[985]/_0_  (.A(\inv_in[985] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[986] ));
 sky130_fd_sc_hd__inv_2 \inv[986]/_0_  (.A(\inv_in[986] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[987] ));
 sky130_fd_sc_hd__inv_2 \inv[987]/_0_  (.A(\inv_in[987] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[988] ));
 sky130_fd_sc_hd__inv_2 \inv[988]/_0_  (.A(\inv_in[988] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[989] ));
 sky130_fd_sc_hd__inv_2 \inv[989]/_0_  (.A(\inv_in[989] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[990] ));
 sky130_fd_sc_hd__inv_2 \inv[98]/_0_  (.A(\inv_in[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[99] ));
 sky130_fd_sc_hd__inv_2 \inv[990]/_0_  (.A(\inv_in[990] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[991] ));
 sky130_fd_sc_hd__inv_2 \inv[991]/_0_  (.A(\inv_in[991] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[992] ));
 sky130_fd_sc_hd__inv_2 \inv[992]/_0_  (.A(\inv_in[992] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[993] ));
 sky130_fd_sc_hd__inv_2 \inv[993]/_0_  (.A(\inv_in[993] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[994] ));
 sky130_fd_sc_hd__inv_2 \inv[994]/_0_  (.A(\inv_in[994] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[995] ));
 sky130_fd_sc_hd__inv_2 \inv[995]/_0_  (.A(\inv_in[995] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[996] ));
 sky130_fd_sc_hd__inv_2 \inv[996]/_0_  (.A(\inv_in[996] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[997] ));
 sky130_fd_sc_hd__inv_2 \inv[997]/_0_  (.A(\inv_in[997] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[998] ));
 sky130_fd_sc_hd__inv_2 \inv[998]/_0_  (.A(\inv_in[998] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[999] ));
 sky130_fd_sc_hd__inv_2 \inv[999]/_0_  (.A(\inv_in[999] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[1000] ));
 sky130_fd_sc_hd__inv_2 \inv[99]/_0_  (.A(\inv_in[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[100] ));
 sky130_fd_sc_hd__inv_2 \inv[9]/_0_  (.A(\inv_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inv_in[10] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__conb_1 tt_um_urish_giant_ringosc_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net3));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[6] = net3;
 assign uio_out[7] = net4;
endmodule
