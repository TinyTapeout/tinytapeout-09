module tt_um_kmakise_sram (clk,
    ena,
    rst_n,
    VDPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VDPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \SRAMController_ins.addr[0] ;
 wire \SRAMController_ins.addr[1] ;
 wire \SRAMController_ins.addr[2] ;
 wire \SRAMController_ins.addr[3] ;
 wire \SRAMController_ins.addr_tmp[0] ;
 wire \SRAMController_ins.addr_tmp[1] ;
 wire \SRAMController_ins.addr_tmp[2] ;
 wire \SRAMController_ins.addr_tmp[3] ;
 wire \SRAMController_ins.csb_n ;
 wire \SRAMController_ins.cur_state[0] ;
 wire \SRAMController_ins.cur_state[1] ;
 wire \SRAMController_ins.cur_state[2] ;
 wire \SRAMController_ins.cur_state[3] ;
 wire \SRAMController_ins.data_tmp[0] ;
 wire \SRAMController_ins.data_tmp[10] ;
 wire \SRAMController_ins.data_tmp[11] ;
 wire \SRAMController_ins.data_tmp[12] ;
 wire \SRAMController_ins.data_tmp[13] ;
 wire \SRAMController_ins.data_tmp[14] ;
 wire \SRAMController_ins.data_tmp[15] ;
 wire \SRAMController_ins.data_tmp[16] ;
 wire \SRAMController_ins.data_tmp[17] ;
 wire \SRAMController_ins.data_tmp[18] ;
 wire \SRAMController_ins.data_tmp[19] ;
 wire \SRAMController_ins.data_tmp[1] ;
 wire \SRAMController_ins.data_tmp[20] ;
 wire \SRAMController_ins.data_tmp[21] ;
 wire \SRAMController_ins.data_tmp[22] ;
 wire \SRAMController_ins.data_tmp[23] ;
 wire \SRAMController_ins.data_tmp[24] ;
 wire \SRAMController_ins.data_tmp[25] ;
 wire \SRAMController_ins.data_tmp[26] ;
 wire \SRAMController_ins.data_tmp[27] ;
 wire \SRAMController_ins.data_tmp[28] ;
 wire \SRAMController_ins.data_tmp[29] ;
 wire \SRAMController_ins.data_tmp[2] ;
 wire \SRAMController_ins.data_tmp[30] ;
 wire \SRAMController_ins.data_tmp[31] ;
 wire \SRAMController_ins.data_tmp[3] ;
 wire \SRAMController_ins.data_tmp[4] ;
 wire \SRAMController_ins.data_tmp[5] ;
 wire \SRAMController_ins.data_tmp[6] ;
 wire \SRAMController_ins.data_tmp[7] ;
 wire \SRAMController_ins.data_tmp[8] ;
 wire \SRAMController_ins.data_tmp[9] ;
 wire \SRAMController_ins.nxt_state[0] ;
 wire \SRAMController_ins.nxt_state[1] ;
 wire \SRAMController_ins.nxt_state[2] ;
 wire \SRAMController_ins.nxt_state[3] ;
 wire \SRAMController_ins.rx_data_out[0] ;
 wire \SRAMController_ins.rx_data_out[1] ;
 wire \SRAMController_ins.rx_data_out[2] ;
 wire \SRAMController_ins.rx_data_out[3] ;
 wire \SRAMController_ins.rx_data_out[4] ;
 wire \SRAMController_ins.rx_data_out[5] ;
 wire \SRAMController_ins.rx_data_out[6] ;
 wire \SRAMController_ins.rx_data_out[7] ;
 wire \SRAMController_ins.rx_valid ;
 wire \SRAMController_ins.sram_addr_from_dpu[0] ;
 wire \SRAMController_ins.sram_addr_from_dpu[1] ;
 wire \SRAMController_ins.sram_addr_from_dpu[2] ;
 wire \SRAMController_ins.sram_addr_from_dpu[3] ;
 wire \SRAMController_ins.sram_data_from_dpu[0] ;
 wire \SRAMController_ins.sram_data_from_dpu[10] ;
 wire \SRAMController_ins.sram_data_from_dpu[11] ;
 wire \SRAMController_ins.sram_data_from_dpu[12] ;
 wire \SRAMController_ins.sram_data_from_dpu[13] ;
 wire \SRAMController_ins.sram_data_from_dpu[14] ;
 wire \SRAMController_ins.sram_data_from_dpu[15] ;
 wire \SRAMController_ins.sram_data_from_dpu[16] ;
 wire \SRAMController_ins.sram_data_from_dpu[17] ;
 wire \SRAMController_ins.sram_data_from_dpu[18] ;
 wire \SRAMController_ins.sram_data_from_dpu[19] ;
 wire \SRAMController_ins.sram_data_from_dpu[1] ;
 wire \SRAMController_ins.sram_data_from_dpu[20] ;
 wire \SRAMController_ins.sram_data_from_dpu[21] ;
 wire \SRAMController_ins.sram_data_from_dpu[22] ;
 wire \SRAMController_ins.sram_data_from_dpu[23] ;
 wire \SRAMController_ins.sram_data_from_dpu[24] ;
 wire \SRAMController_ins.sram_data_from_dpu[25] ;
 wire \SRAMController_ins.sram_data_from_dpu[26] ;
 wire \SRAMController_ins.sram_data_from_dpu[27] ;
 wire \SRAMController_ins.sram_data_from_dpu[28] ;
 wire \SRAMController_ins.sram_data_from_dpu[29] ;
 wire \SRAMController_ins.sram_data_from_dpu[2] ;
 wire \SRAMController_ins.sram_data_from_dpu[30] ;
 wire \SRAMController_ins.sram_data_from_dpu[31] ;
 wire \SRAMController_ins.sram_data_from_dpu[3] ;
 wire \SRAMController_ins.sram_data_from_dpu[4] ;
 wire \SRAMController_ins.sram_data_from_dpu[5] ;
 wire \SRAMController_ins.sram_data_from_dpu[6] ;
 wire \SRAMController_ins.sram_data_from_dpu[7] ;
 wire \SRAMController_ins.sram_data_from_dpu[8] ;
 wire \SRAMController_ins.sram_data_from_dpu[9] ;
 wire \SRAMController_ins.sram_data_in[0] ;
 wire \SRAMController_ins.sram_data_in[10] ;
 wire \SRAMController_ins.sram_data_in[11] ;
 wire \SRAMController_ins.sram_data_in[12] ;
 wire \SRAMController_ins.sram_data_in[13] ;
 wire \SRAMController_ins.sram_data_in[14] ;
 wire \SRAMController_ins.sram_data_in[15] ;
 wire \SRAMController_ins.sram_data_in[16] ;
 wire \SRAMController_ins.sram_data_in[17] ;
 wire \SRAMController_ins.sram_data_in[18] ;
 wire \SRAMController_ins.sram_data_in[19] ;
 wire \SRAMController_ins.sram_data_in[1] ;
 wire \SRAMController_ins.sram_data_in[20] ;
 wire \SRAMController_ins.sram_data_in[21] ;
 wire \SRAMController_ins.sram_data_in[22] ;
 wire \SRAMController_ins.sram_data_in[23] ;
 wire \SRAMController_ins.sram_data_in[24] ;
 wire \SRAMController_ins.sram_data_in[25] ;
 wire \SRAMController_ins.sram_data_in[26] ;
 wire \SRAMController_ins.sram_data_in[27] ;
 wire \SRAMController_ins.sram_data_in[28] ;
 wire \SRAMController_ins.sram_data_in[29] ;
 wire \SRAMController_ins.sram_data_in[2] ;
 wire \SRAMController_ins.sram_data_in[30] ;
 wire \SRAMController_ins.sram_data_in[31] ;
 wire \SRAMController_ins.sram_data_in[3] ;
 wire \SRAMController_ins.sram_data_in[4] ;
 wire \SRAMController_ins.sram_data_in[5] ;
 wire \SRAMController_ins.sram_data_in[6] ;
 wire \SRAMController_ins.sram_data_in[7] ;
 wire \SRAMController_ins.sram_data_in[8] ;
 wire \SRAMController_ins.sram_data_in[9] ;
 wire \SRAMController_ins.sram_data_out[0] ;
 wire \SRAMController_ins.sram_data_out[10] ;
 wire \SRAMController_ins.sram_data_out[11] ;
 wire \SRAMController_ins.sram_data_out[12] ;
 wire \SRAMController_ins.sram_data_out[13] ;
 wire \SRAMController_ins.sram_data_out[14] ;
 wire \SRAMController_ins.sram_data_out[15] ;
 wire \SRAMController_ins.sram_data_out[16] ;
 wire \SRAMController_ins.sram_data_out[17] ;
 wire \SRAMController_ins.sram_data_out[18] ;
 wire \SRAMController_ins.sram_data_out[19] ;
 wire \SRAMController_ins.sram_data_out[1] ;
 wire \SRAMController_ins.sram_data_out[20] ;
 wire \SRAMController_ins.sram_data_out[21] ;
 wire \SRAMController_ins.sram_data_out[22] ;
 wire \SRAMController_ins.sram_data_out[23] ;
 wire \SRAMController_ins.sram_data_out[24] ;
 wire \SRAMController_ins.sram_data_out[25] ;
 wire \SRAMController_ins.sram_data_out[26] ;
 wire \SRAMController_ins.sram_data_out[27] ;
 wire \SRAMController_ins.sram_data_out[28] ;
 wire \SRAMController_ins.sram_data_out[29] ;
 wire \SRAMController_ins.sram_data_out[2] ;
 wire \SRAMController_ins.sram_data_out[30] ;
 wire \SRAMController_ins.sram_data_out[31] ;
 wire \SRAMController_ins.sram_data_out[3] ;
 wire \SRAMController_ins.sram_data_out[4] ;
 wire \SRAMController_ins.sram_data_out[5] ;
 wire \SRAMController_ins.sram_data_out[6] ;
 wire \SRAMController_ins.sram_data_out[7] ;
 wire \SRAMController_ins.sram_data_out[8] ;
 wire \SRAMController_ins.sram_data_out[9] ;
 wire \SRAMController_ins.sram_tmp[0] ;
 wire \SRAMController_ins.sram_tmp[10] ;
 wire \SRAMController_ins.sram_tmp[11] ;
 wire \SRAMController_ins.sram_tmp[12] ;
 wire \SRAMController_ins.sram_tmp[13] ;
 wire \SRAMController_ins.sram_tmp[14] ;
 wire \SRAMController_ins.sram_tmp[15] ;
 wire \SRAMController_ins.sram_tmp[16] ;
 wire \SRAMController_ins.sram_tmp[17] ;
 wire \SRAMController_ins.sram_tmp[18] ;
 wire \SRAMController_ins.sram_tmp[19] ;
 wire \SRAMController_ins.sram_tmp[1] ;
 wire \SRAMController_ins.sram_tmp[20] ;
 wire \SRAMController_ins.sram_tmp[21] ;
 wire \SRAMController_ins.sram_tmp[22] ;
 wire \SRAMController_ins.sram_tmp[23] ;
 wire \SRAMController_ins.sram_tmp[24] ;
 wire \SRAMController_ins.sram_tmp[25] ;
 wire \SRAMController_ins.sram_tmp[26] ;
 wire \SRAMController_ins.sram_tmp[27] ;
 wire \SRAMController_ins.sram_tmp[28] ;
 wire \SRAMController_ins.sram_tmp[29] ;
 wire \SRAMController_ins.sram_tmp[2] ;
 wire \SRAMController_ins.sram_tmp[30] ;
 wire \SRAMController_ins.sram_tmp[31] ;
 wire \SRAMController_ins.sram_tmp[3] ;
 wire \SRAMController_ins.sram_tmp[4] ;
 wire \SRAMController_ins.sram_tmp[5] ;
 wire \SRAMController_ins.sram_tmp[6] ;
 wire \SRAMController_ins.sram_tmp[7] ;
 wire \SRAMController_ins.sram_tmp[8] ;
 wire \SRAMController_ins.sram_tmp[9] ;
 wire \SRAMController_ins.tx_ready ;
 wire \SRAMController_ins.uart_ready ;
 wire \SRAMController_ins.we_n ;
 wire \UARTReceiver_ins.bitIndex[0] ;
 wire \UARTReceiver_ins.bitIndex[1] ;
 wire \UARTReceiver_ins.bitIndex[2] ;
 wire \UARTReceiver_ins.data[0] ;
 wire \UARTReceiver_ins.data[1] ;
 wire \UARTReceiver_ins.data[2] ;
 wire \UARTReceiver_ins.data[3] ;
 wire \UARTReceiver_ins.data[4] ;
 wire \UARTReceiver_ins.data[5] ;
 wire \UARTReceiver_ins.data[6] ;
 wire \UARTReceiver_ins.data[7] ;
 wire \UARTReceiver_ins.error ;
 wire \UARTReceiver_ins.inputReg[0] ;
 wire \UARTReceiver_ins.inputReg[1] ;
 wire \UARTReceiver_ins.inputReg[2] ;
 wire \UARTReceiver_ins.out_latched ;
 wire \UARTReceiver_ins.overrun ;
 wire \UARTReceiver_ins.rxCounter[0] ;
 wire \UARTReceiver_ins.rxCounter[1] ;
 wire \UARTReceiver_ins.rxCounter[2] ;
 wire \UARTReceiver_ins.rxCounter[3] ;
 wire \UARTReceiver_ins.rxCounter[4] ;
 wire \UARTReceiver_ins.rxCounter[5] ;
 wire \UARTReceiver_ins.rxCounter[6] ;
 wire \UARTReceiver_ins.rxCounter[7] ;
 wire \UARTReceiver_ins.sampleCount[0] ;
 wire \UARTReceiver_ins.sampleCount[1] ;
 wire \UARTReceiver_ins.sampleCount[2] ;
 wire \UARTReceiver_ins.sampleCount[3] ;
 wire \UARTReceiver_ins.state[0] ;
 wire \UARTReceiver_ins.state[1] ;
 wire \UARTReceiver_ins.state[2] ;
 wire \UARTReceiver_ins.state[3] ;
 wire \UARTTransmitter_ins.bitIndex[0] ;
 wire \UARTTransmitter_ins.bitIndex[1] ;
 wire \UARTTransmitter_ins.bitIndex[2] ;
 wire \UARTTransmitter_ins.data[0] ;
 wire \UARTTransmitter_ins.data[1] ;
 wire \UARTTransmitter_ins.data[2] ;
 wire \UARTTransmitter_ins.data[3] ;
 wire \UARTTransmitter_ins.data[4] ;
 wire \UARTTransmitter_ins.data[5] ;
 wire \UARTTransmitter_ins.data[6] ;
 wire \UARTTransmitter_ins.data[7] ;
 wire \UARTTransmitter_ins.out ;
 wire \UARTTransmitter_ins.state[0] ;
 wire \UARTTransmitter_ins.state[1] ;
 wire \UARTTransmitter_ins.state[2] ;
 wire \UARTTransmitter_ins.state[3] ;
 wire \UARTTransmitter_ins.txCounter[0] ;
 wire \UARTTransmitter_ins.txCounter[10] ;
 wire \UARTTransmitter_ins.txCounter[11] ;
 wire \UARTTransmitter_ins.txCounter[1] ;
 wire \UARTTransmitter_ins.txCounter[2] ;
 wire \UARTTransmitter_ins.txCounter[3] ;
 wire \UARTTransmitter_ins.txCounter[4] ;
 wire \UARTTransmitter_ins.txCounter[5] ;
 wire \UARTTransmitter_ins.txCounter[6] ;
 wire \UARTTransmitter_ins.txCounter[7] ;
 wire \UARTTransmitter_ins.txCounter[8] ;
 wire \UARTTransmitter_ins.txCounter[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire net67;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire \dpu_ins.cur_cmd[5] ;
 wire \dpu_ins.cur_cmd[6] ;
 wire \dpu_ins.cur_state[0] ;
 wire \dpu_ins.cur_state[1] ;
 wire \dpu_ins.data_in[0] ;
 wire \dpu_ins.data_in[10] ;
 wire \dpu_ins.data_in[11] ;
 wire \dpu_ins.data_in[12] ;
 wire \dpu_ins.data_in[13] ;
 wire \dpu_ins.data_in[14] ;
 wire \dpu_ins.data_in[15] ;
 wire \dpu_ins.data_in[16] ;
 wire \dpu_ins.data_in[17] ;
 wire \dpu_ins.data_in[18] ;
 wire \dpu_ins.data_in[19] ;
 wire \dpu_ins.data_in[1] ;
 wire \dpu_ins.data_in[20] ;
 wire \dpu_ins.data_in[21] ;
 wire \dpu_ins.data_in[22] ;
 wire \dpu_ins.data_in[23] ;
 wire \dpu_ins.data_in[24] ;
 wire \dpu_ins.data_in[25] ;
 wire \dpu_ins.data_in[26] ;
 wire \dpu_ins.data_in[27] ;
 wire \dpu_ins.data_in[28] ;
 wire \dpu_ins.data_in[29] ;
 wire \dpu_ins.data_in[2] ;
 wire \dpu_ins.data_in[30] ;
 wire \dpu_ins.data_in[31] ;
 wire \dpu_ins.data_in[3] ;
 wire \dpu_ins.data_in[4] ;
 wire \dpu_ins.data_in[5] ;
 wire \dpu_ins.data_in[6] ;
 wire \dpu_ins.data_in[7] ;
 wire \dpu_ins.data_in[8] ;
 wire \dpu_ins.data_in[9] ;
 wire \dpu_ins.data_out[0] ;
 wire \dpu_ins.data_out[10] ;
 wire \dpu_ins.data_out[11] ;
 wire \dpu_ins.data_out[12] ;
 wire \dpu_ins.data_out[13] ;
 wire \dpu_ins.data_out[14] ;
 wire \dpu_ins.data_out[15] ;
 wire \dpu_ins.data_out[16] ;
 wire \dpu_ins.data_out[17] ;
 wire \dpu_ins.data_out[18] ;
 wire \dpu_ins.data_out[19] ;
 wire \dpu_ins.data_out[1] ;
 wire \dpu_ins.data_out[20] ;
 wire \dpu_ins.data_out[21] ;
 wire \dpu_ins.data_out[22] ;
 wire \dpu_ins.data_out[23] ;
 wire \dpu_ins.data_out[24] ;
 wire \dpu_ins.data_out[25] ;
 wire \dpu_ins.data_out[26] ;
 wire \dpu_ins.data_out[27] ;
 wire \dpu_ins.data_out[28] ;
 wire \dpu_ins.data_out[29] ;
 wire \dpu_ins.data_out[2] ;
 wire \dpu_ins.data_out[30] ;
 wire \dpu_ins.data_out[31] ;
 wire \dpu_ins.data_out[3] ;
 wire \dpu_ins.data_out[4] ;
 wire \dpu_ins.data_out[5] ;
 wire \dpu_ins.data_out[6] ;
 wire \dpu_ins.data_out[7] ;
 wire \dpu_ins.data_out[8] ;
 wire \dpu_ins.data_out[9] ;
 wire \dpu_ins.nxt_state[0] ;
 wire \dpu_ins.nxt_state[1] ;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire clknet_leaf_0_clk;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;

 sky130_fd_sc_hd__or2_1 _0787_ (.A(\UARTReceiver_ins.rxCounter[0] ),
    .B(\UARTReceiver_ins.rxCounter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0382_));
 sky130_fd_sc_hd__o41a_1 _0788_ (.A1(\UARTReceiver_ins.rxCounter[4] ),
    .A2(\UARTReceiver_ins.rxCounter[3] ),
    .A3(\UARTReceiver_ins.rxCounter[2] ),
    .A4(_0382_),
    .B1(\UARTReceiver_ins.rxCounter[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0383_));
 sky130_fd_sc_hd__o21a_2 _0789_ (.A1(\UARTReceiver_ins.rxCounter[6] ),
    .A2(_0383_),
    .B1(\UARTReceiver_ins.rxCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0384_));
 sky130_fd_sc_hd__and2_1 _0790_ (.A(\UARTReceiver_ins.inputReg[1] ),
    .B(\UARTReceiver_ins.inputReg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0385_));
 sky130_fd_sc_hd__nand2_1 _0791_ (.A(\UARTReceiver_ins.inputReg[2] ),
    .B(_0385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0386_));
 sky130_fd_sc_hd__and4_2 _0792_ (.A(\UARTReceiver_ins.sampleCount[3] ),
    .B(\UARTReceiver_ins.sampleCount[2] ),
    .C(\UARTReceiver_ins.sampleCount[1] ),
    .D(\UARTReceiver_ins.sampleCount[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0387_));
 sky130_fd_sc_hd__o21ai_4 _0793_ (.A1(\UARTReceiver_ins.rxCounter[6] ),
    .A2(_0383_),
    .B1(\UARTReceiver_ins.rxCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0388_));
 sky130_fd_sc_hd__nand2_2 _0794_ (.A(net25),
    .B(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0389_));
 sky130_fd_sc_hd__nand2_2 _0795_ (.A(net25),
    .B(_0384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0390_));
 sky130_fd_sc_hd__or2_1 _0796_ (.A(\UARTReceiver_ins.sampleCount[1] ),
    .B(\UARTReceiver_ins.sampleCount[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0391_));
 sky130_fd_sc_hd__a21oi_1 _0797_ (.A1(\UARTReceiver_ins.sampleCount[2] ),
    .A2(_0391_),
    .B1(\UARTReceiver_ins.sampleCount[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0392_));
 sky130_fd_sc_hd__or3_1 _0798_ (.A(\UARTReceiver_ins.sampleCount[3] ),
    .B(\UARTReceiver_ins.sampleCount[2] ),
    .C(_0391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0393_));
 sky130_fd_sc_hd__or3_1 _0799_ (.A(\UARTReceiver_ins.inputReg[2] ),
    .B(\UARTReceiver_ins.inputReg[1] ),
    .C(\UARTReceiver_ins.inputReg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0394_));
 sky130_fd_sc_hd__and4_1 _0800_ (.A(\UARTReceiver_ins.state[2] ),
    .B(_0392_),
    .C(_0393_),
    .D(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0395_));
 sky130_fd_sc_hd__o22a_1 _0801_ (.A1(net16),
    .A2(_0389_),
    .B1(_0390_),
    .B2(_0395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0396_));
 sky130_fd_sc_hd__a41o_1 _0802_ (.A1(net14),
    .A2(_0384_),
    .A3(_0386_),
    .A4(_0387_),
    .B1(_0396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0000_));
 sky130_fd_sc_hd__inv_2 _0803_ (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0397_));
 sky130_fd_sc_hd__clkbuf_4 _0804_ (.A(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0398_));
 sky130_fd_sc_hd__inv_2 _0805_ (.A(\UARTReceiver_ins.state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0399_));
 sky130_fd_sc_hd__nand3_1 _0806_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .B(net19),
    .C(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0400_));
 sky130_fd_sc_hd__nand2_1 _0807_ (.A(_0384_),
    .B(_0387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0401_));
 sky130_fd_sc_hd__nor2_1 _0808_ (.A(_0400_),
    .B(_0401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _0809_ (.A(\UARTReceiver_ins.state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0403_));
 sky130_fd_sc_hd__or3_1 _0810_ (.A(_0403_),
    .B(_0390_),
    .C(_0392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0404_));
 sky130_fd_sc_hd__o31ai_1 _0811_ (.A1(_0398_),
    .A2(_0399_),
    .A3(_0402_),
    .B1(_0404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0001_));
 sky130_fd_sc_hd__a21o_1 _0812_ (.A1(\UARTTransmitter_ins.txCounter[1] ),
    .A2(\UARTTransmitter_ins.txCounter[0] ),
    .B1(\UARTTransmitter_ins.txCounter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0405_));
 sky130_fd_sc_hd__a21o_1 _0813_ (.A1(\UARTTransmitter_ins.txCounter[3] ),
    .A2(_0405_),
    .B1(\UARTTransmitter_ins.txCounter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0406_));
 sky130_fd_sc_hd__a2111o_1 _0814_ (.A1(\UARTTransmitter_ins.txCounter[5] ),
    .A2(_0406_),
    .B1(\UARTTransmitter_ins.txCounter[8] ),
    .C1(\UARTTransmitter_ins.txCounter[7] ),
    .D1(\UARTTransmitter_ins.txCounter[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0407_));
 sky130_fd_sc_hd__a21o_1 _0815_ (.A1(\UARTTransmitter_ins.txCounter[9] ),
    .A2(_0407_),
    .B1(\UARTTransmitter_ins.txCounter[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0408_));
 sky130_fd_sc_hd__and2_2 _0816_ (.A(\UARTTransmitter_ins.txCounter[11] ),
    .B(_0408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0409_));
 sky130_fd_sc_hd__inv_2 _0817_ (.A(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0410_));
 sky130_fd_sc_hd__or2_2 _0818_ (.A(\SRAMController_ins.cur_state[2] ),
    .B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0411_));
 sky130_fd_sc_hd__nand2b_4 _0819_ (.A_N(\SRAMController_ins.cur_state[0] ),
    .B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0412_));
 sky130_fd_sc_hd__nor2_4 _0820_ (.A(_0411_),
    .B(_0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0413_));
 sky130_fd_sc_hd__or2b_1 _0821_ (.A(\SRAMController_ins.cur_state[0] ),
    .B_N(\SRAMController_ins.cur_state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0414_));
 sky130_fd_sc_hd__nor2_1 _0822_ (.A(\SRAMController_ins.cur_state[3] ),
    .B(_0414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0415_));
 sky130_fd_sc_hd__and2b_1 _0823_ (.A_N(net9),
    .B(_0415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0416_));
 sky130_fd_sc_hd__nand2_1 _0824_ (.A(net9),
    .B(\SRAMController_ins.cur_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0417_));
 sky130_fd_sc_hd__nor2_1 _0825_ (.A(_0411_),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0418_));
 sky130_fd_sc_hd__nand2_1 _0826_ (.A(\SRAMController_ins.cur_state[0] ),
    .B(\SRAMController_ins.cur_state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0419_));
 sky130_fd_sc_hd__nor2_1 _0827_ (.A(net7),
    .B(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0420_));
 sky130_fd_sc_hd__nor2b_4 _0828_ (.A(net9),
    .B_N(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0421_));
 sky130_fd_sc_hd__or4_1 _0829_ (.A(_0413_),
    .B(_0416_),
    .C(_0418_),
    .D(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_2 _0830_ (.A(net17),
    .B(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_2 _0831_ (.A(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0424_));
 sky130_fd_sc_hd__nor2_1 _0832_ (.A(_0397_),
    .B(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0425_));
 sky130_fd_sc_hd__and2_1 _0833_ (.A(\UARTTransmitter_ins.bitIndex[1] ),
    .B(\UARTTransmitter_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0426_));
 sky130_fd_sc_hd__and4_1 _0834_ (.A(\UARTTransmitter_ins.bitIndex[2] ),
    .B(_0409_),
    .C(_0426_),
    .D(_0425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0427_));
 sky130_fd_sc_hd__a32o_1 _0835_ (.A1(net88),
    .A2(_0410_),
    .A3(_0425_),
    .B1(_0427_),
    .B2(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_2 _0836_ (.A(_0410_),
    .B(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0428_));
 sky130_fd_sc_hd__nor2_1 _0837_ (.A(_0397_),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0429_));
 sky130_fd_sc_hd__clkbuf_2 _0838_ (.A(_0429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0430_));
 sky130_fd_sc_hd__o21a_1 _0839_ (.A1(net68),
    .A2(_0424_),
    .B1(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _0840_ (.A(\UARTTransmitter_ins.bitIndex[2] ),
    .B(_0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0431_));
 sky130_fd_sc_hd__o211a_1 _0841_ (.A1(_0410_),
    .A2(_0431_),
    .B1(_0425_),
    .C1(\UARTTransmitter_ins.state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0432_));
 sky130_fd_sc_hd__a31o_1 _0842_ (.A1(net28),
    .A2(net68),
    .A3(_0428_),
    .B1(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0005_));
 sky130_fd_sc_hd__a221o_1 _0843_ (.A1(\UARTTransmitter_ins.state[0] ),
    .A2(_0423_),
    .B1(_0428_),
    .B2(net88),
    .C1(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0004_));
 sky130_fd_sc_hd__and3_1 _0844_ (.A(net14),
    .B(net25),
    .C(_0401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0433_));
 sky130_fd_sc_hd__a31o_1 _0845_ (.A1(net25),
    .A2(net15),
    .A3(_0402_),
    .B1(_0433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0003_));
 sky130_fd_sc_hd__nor2_2 _0846_ (.A(_0397_),
    .B(_0384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0434_));
 sky130_fd_sc_hd__nand2_1 _0847_ (.A(\UARTReceiver_ins.state[2] ),
    .B(_0392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0435_));
 sky130_fd_sc_hd__nor2_1 _0848_ (.A(_0394_),
    .B(_0435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0436_));
 sky130_fd_sc_hd__and4_1 _0849_ (.A(net14),
    .B(\UARTReceiver_ins.inputReg[2] ),
    .C(_0385_),
    .D(_0387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0437_));
 sky130_fd_sc_hd__nor3b_1 _0850_ (.A(_0403_),
    .B(_0393_),
    .C_N(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0438_));
 sky130_fd_sc_hd__or2_1 _0851_ (.A(_0437_),
    .B(_0438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0439_));
 sky130_fd_sc_hd__o21ba_1 _0852_ (.A1(net16),
    .A2(_0439_),
    .B1_N(_0390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0440_));
 sky130_fd_sc_hd__a221o_1 _0853_ (.A1(\UARTReceiver_ins.state[2] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(net25),
    .C1(_0440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0002_));
 sky130_fd_sc_hd__nor2_1 _0854_ (.A(\SRAMController_ins.cur_state[2] ),
    .B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0441_));
 sky130_fd_sc_hd__nor2_1 _0855_ (.A(net8),
    .B(\SRAMController_ins.cur_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0442_));
 sky130_fd_sc_hd__and2_1 _0856_ (.A(_0441_),
    .B(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0443_));
 sky130_fd_sc_hd__buf_1 _0857_ (.A(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.uart_ready ));
 sky130_fd_sc_hd__and2_1 _0858_ (.A(net10),
    .B(\dpu_ins.cur_cmd[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0444_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0859_ (.A(_0444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_4 _0860_ (.A(_0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0446_));
 sky130_fd_sc_hd__a2bb2o_1 _0861_ (.A1_N(\dpu_ins.data_in[0] ),
    .A2_N(net10),
    .B1(\dpu_ins.data_in[1] ),
    .B2(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[0] ));
 sky130_fd_sc_hd__inv_2 _0862_ (.A(_0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0447_));
 sky130_fd_sc_hd__and2b_1 _0863_ (.A_N(net10),
    .B(\dpu_ins.cur_cmd[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_2 _0864_ (.A(_0448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0449_));
 sky130_fd_sc_hd__buf_2 _0865_ (.A(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_4 _0866_ (.A(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_4 _0867_ (.A(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_4 _0868_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0453_));
 sky130_fd_sc_hd__buf_2 _0869_ (.A(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0454_));
 sky130_fd_sc_hd__buf_4 _0870_ (.A(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0455_));
 sky130_fd_sc_hd__and2_1 _0871_ (.A(\dpu_ins.data_in[1] ),
    .B(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0456_));
 sky130_fd_sc_hd__nor2_1 _0872_ (.A(\dpu_ins.data_in[1] ),
    .B(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0457_));
 sky130_fd_sc_hd__or3_1 _0873_ (.A(net10),
    .B(_0456_),
    .C(_0457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0458_));
 sky130_fd_sc_hd__a2bb2o_1 _0874_ (.A1_N(\dpu_ins.data_in[0] ),
    .A2_N(_0458_),
    .B1(_0445_),
    .B2(\dpu_ins.data_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0459_));
 sky130_fd_sc_hd__a31o_1 _0875_ (.A1(\dpu_ins.data_in[0] ),
    .A2(_0447_),
    .A3(_0458_),
    .B1(_0459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[1] ));
 sky130_fd_sc_hd__inv_2 _0876_ (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0460_));
 sky130_fd_sc_hd__nor2_1 _0877_ (.A(_0460_),
    .B(\dpu_ins.cur_cmd[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0461_));
 sky130_fd_sc_hd__buf_4 _0878_ (.A(_0461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0462_));
 sky130_fd_sc_hd__xnor2_1 _0879_ (.A(\dpu_ins.data_in[2] ),
    .B(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0463_));
 sky130_fd_sc_hd__a21oi_1 _0880_ (.A1(\dpu_ins.data_in[1] ),
    .A2(_0449_),
    .B1(\dpu_ins.data_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0464_));
 sky130_fd_sc_hd__nor3_1 _0881_ (.A(_0457_),
    .B(_0463_),
    .C(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0465_));
 sky130_fd_sc_hd__o21a_1 _0882_ (.A1(_0457_),
    .A2(_0464_),
    .B1(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0466_));
 sky130_fd_sc_hd__nor3_1 _0883_ (.A(net10),
    .B(_0465_),
    .C(_0466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0467_));
 sky130_fd_sc_hd__a221o_1 _0884_ (.A1(\dpu_ins.data_in[3] ),
    .A2(_0446_),
    .B1(_0462_),
    .B2(\dpu_ins.data_in[1] ),
    .C1(_0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[2] ));
 sky130_fd_sc_hd__a21o_1 _0885_ (.A1(\dpu_ins.data_in[2] ),
    .A2(_0455_),
    .B1(_0465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0468_));
 sky130_fd_sc_hd__xor2_1 _0886_ (.A(\dpu_ins.data_in[3] ),
    .B(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0469_));
 sky130_fd_sc_hd__buf_4 _0887_ (.A(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0470_));
 sky130_fd_sc_hd__o21a_1 _0888_ (.A1(_0468_),
    .A2(_0469_),
    .B1(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0471_));
 sky130_fd_sc_hd__a21boi_1 _0889_ (.A1(_0468_),
    .A2(_0469_),
    .B1_N(_0471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0472_));
 sky130_fd_sc_hd__a221o_1 _0890_ (.A1(\dpu_ins.data_in[4] ),
    .A2(_0446_),
    .B1(_0462_),
    .B2(\dpu_ins.data_in[2] ),
    .C1(_0472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[3] ));
 sky130_fd_sc_hd__clkbuf_4 _0891_ (.A(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_1 _0892_ (.A(\dpu_ins.data_in[2] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_1 _0893_ (.A(\dpu_ins.data_in[3] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0475_));
 sky130_fd_sc_hd__or4b_1 _0894_ (.A(_0457_),
    .B(_0463_),
    .C(_0464_),
    .D_N(_0469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_1 _0895_ (.A(\dpu_ins.data_in[4] ),
    .B(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0477_));
 sky130_fd_sc_hd__or2_1 _0896_ (.A(\dpu_ins.data_in[4] ),
    .B(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0478_));
 sky130_fd_sc_hd__nand2_1 _0897_ (.A(_0477_),
    .B(_0478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0479_));
 sky130_fd_sc_hd__a31o_1 _0898_ (.A1(_0474_),
    .A2(_0475_),
    .A3(_0476_),
    .B1(_0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0480_));
 sky130_fd_sc_hd__a41oi_1 _0899_ (.A1(_0474_),
    .A2(_0475_),
    .A3(_0479_),
    .A4(_0476_),
    .B1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0481_));
 sky130_fd_sc_hd__buf_4 _0900_ (.A(_0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0482_));
 sky130_fd_sc_hd__buf_4 _0901_ (.A(_0461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0483_));
 sky130_fd_sc_hd__a22o_1 _0902_ (.A1(\dpu_ins.data_in[5] ),
    .A2(_0482_),
    .B1(_0483_),
    .B2(\dpu_ins.data_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0484_));
 sky130_fd_sc_hd__a21o_1 _0903_ (.A1(_0480_),
    .A2(_0481_),
    .B1(_0484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[4] ));
 sky130_fd_sc_hd__and2_1 _0904_ (.A(\dpu_ins.data_in[5] ),
    .B(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0485_));
 sky130_fd_sc_hd__nor2_1 _0905_ (.A(\dpu_ins.data_in[5] ),
    .B(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0486_));
 sky130_fd_sc_hd__or2_1 _0906_ (.A(_0485_),
    .B(_0486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0487_));
 sky130_fd_sc_hd__a21oi_1 _0907_ (.A1(_0477_),
    .A2(_0480_),
    .B1(_0487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0488_));
 sky130_fd_sc_hd__a31o_1 _0908_ (.A1(_0477_),
    .A2(_0480_),
    .A3(_0487_),
    .B1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0489_));
 sky130_fd_sc_hd__nor2_1 _0909_ (.A(_0488_),
    .B(_0489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0490_));
 sky130_fd_sc_hd__a221o_1 _0910_ (.A1(\dpu_ins.data_in[6] ),
    .A2(_0446_),
    .B1(_0462_),
    .B2(\dpu_ins.data_in[4] ),
    .C1(_0490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[5] ));
 sky130_fd_sc_hd__nand2_1 _0911_ (.A(\dpu_ins.data_in[6] ),
    .B(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0491_));
 sky130_fd_sc_hd__or2_1 _0912_ (.A(\dpu_ins.data_in[6] ),
    .B(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_1 _0913_ (.A(_0491_),
    .B(_0492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0493_));
 sky130_fd_sc_hd__o21ai_1 _0914_ (.A1(\dpu_ins.data_in[4] ),
    .A2(\dpu_ins.data_in[5] ),
    .B1(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0494_));
 sky130_fd_sc_hd__a21o_1 _0915_ (.A1(_0480_),
    .A2(_0494_),
    .B1(_0486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0495_));
 sky130_fd_sc_hd__or2_1 _0916_ (.A(_0493_),
    .B(_0495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0496_));
 sky130_fd_sc_hd__nand2_1 _0917_ (.A(_0493_),
    .B(_0495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0497_));
 sky130_fd_sc_hd__a22o_1 _0918_ (.A1(\dpu_ins.data_in[7] ),
    .A2(_0482_),
    .B1(_0483_),
    .B2(\dpu_ins.data_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0498_));
 sky130_fd_sc_hd__a31o_1 _0919_ (.A1(_0470_),
    .A2(_0496_),
    .A3(_0497_),
    .B1(_0498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[6] ));
 sky130_fd_sc_hd__xnor2_1 _0920_ (.A(\dpu_ins.data_in[7] ),
    .B(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0499_));
 sky130_fd_sc_hd__a21oi_1 _0921_ (.A1(_0491_),
    .A2(_0496_),
    .B1(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0500_));
 sky130_fd_sc_hd__a31o_1 _0922_ (.A1(_0491_),
    .A2(_0496_),
    .A3(_0499_),
    .B1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0501_));
 sky130_fd_sc_hd__nor2_1 _0923_ (.A(_0500_),
    .B(_0501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0502_));
 sky130_fd_sc_hd__a221o_1 _0924_ (.A1(\dpu_ins.data_in[8] ),
    .A2(_0446_),
    .B1(_0462_),
    .B2(\dpu_ins.data_in[6] ),
    .C1(_0502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[7] ));
 sky130_fd_sc_hd__or3_1 _0925_ (.A(_0487_),
    .B(_0493_),
    .C(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0503_));
 sky130_fd_sc_hd__o21ai_1 _0926_ (.A1(\dpu_ins.data_in[6] ),
    .A2(\dpu_ins.data_in[7] ),
    .B1(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0504_));
 sky130_fd_sc_hd__o211a_1 _0927_ (.A1(_0480_),
    .A2(_0503_),
    .B1(_0504_),
    .C1(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0505_));
 sky130_fd_sc_hd__nand2_1 _0928_ (.A(\dpu_ins.data_in[8] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0506_));
 sky130_fd_sc_hd__or2_1 _0929_ (.A(\dpu_ins.data_in[8] ),
    .B(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0507_));
 sky130_fd_sc_hd__nand2_1 _0930_ (.A(_0506_),
    .B(_0507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0508_));
 sky130_fd_sc_hd__or2_1 _0931_ (.A(_0505_),
    .B(_0508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_1 _0932_ (.A(_0505_),
    .B(_0508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0510_));
 sky130_fd_sc_hd__a22o_1 _0933_ (.A1(\dpu_ins.data_in[9] ),
    .A2(_0482_),
    .B1(_0483_),
    .B2(\dpu_ins.data_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0511_));
 sky130_fd_sc_hd__a31o_1 _0934_ (.A1(_0470_),
    .A2(_0509_),
    .A3(_0510_),
    .B1(_0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[8] ));
 sky130_fd_sc_hd__o21ai_1 _0935_ (.A1(_0505_),
    .A2(_0508_),
    .B1(_0506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0512_));
 sky130_fd_sc_hd__or2_1 _0936_ (.A(\dpu_ins.data_in[9] ),
    .B(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _0937_ (.A(\dpu_ins.data_in[9] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0514_));
 sky130_fd_sc_hd__nand2_1 _0938_ (.A(_0513_),
    .B(_0514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0515_));
 sky130_fd_sc_hd__xor2_1 _0939_ (.A(_0512_),
    .B(_0515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0516_));
 sky130_fd_sc_hd__nor2_1 _0940_ (.A(net11),
    .B(_0516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0517_));
 sky130_fd_sc_hd__a221o_1 _0941_ (.A1(\dpu_ins.data_in[10] ),
    .A2(_0446_),
    .B1(_0462_),
    .B2(\dpu_ins.data_in[8] ),
    .C1(_0517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[9] ));
 sky130_fd_sc_hd__nand2_1 _0942_ (.A(\dpu_ins.data_in[10] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0518_));
 sky130_fd_sc_hd__or2_1 _0943_ (.A(\dpu_ins.data_in[10] ),
    .B(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0519_));
 sky130_fd_sc_hd__nand2_1 _0944_ (.A(_0518_),
    .B(_0519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0520_));
 sky130_fd_sc_hd__and2_1 _0945_ (.A(\dpu_ins.data_in[9] ),
    .B(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0521_));
 sky130_fd_sc_hd__a21oi_1 _0946_ (.A1(_0512_),
    .A2(_0513_),
    .B1(_0521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0522_));
 sky130_fd_sc_hd__a21oi_1 _0947_ (.A1(_0520_),
    .A2(_0522_),
    .B1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0523_));
 sky130_fd_sc_hd__o21a_1 _0948_ (.A1(_0520_),
    .A2(_0522_),
    .B1(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0524_));
 sky130_fd_sc_hd__a221o_1 _0949_ (.A1(\dpu_ins.data_in[11] ),
    .A2(_0446_),
    .B1(_0462_),
    .B2(\dpu_ins.data_in[9] ),
    .C1(_0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[10] ));
 sky130_fd_sc_hd__xnor2_1 _0950_ (.A(\dpu_ins.data_in[11] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0525_));
 sky130_fd_sc_hd__o21ai_1 _0951_ (.A1(_0520_),
    .A2(_0522_),
    .B1(_0518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0526_));
 sky130_fd_sc_hd__xor2_1 _0952_ (.A(_0525_),
    .B(_0526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0527_));
 sky130_fd_sc_hd__nor2_1 _0953_ (.A(net11),
    .B(_0527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0528_));
 sky130_fd_sc_hd__a221o_1 _0954_ (.A1(\dpu_ins.data_in[12] ),
    .A2(_0446_),
    .B1(_0462_),
    .B2(\dpu_ins.data_in[10] ),
    .C1(_0528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[11] ));
 sky130_fd_sc_hd__and2_1 _0955_ (.A(\dpu_ins.data_in[12] ),
    .B(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0529_));
 sky130_fd_sc_hd__nor2_1 _0956_ (.A(\dpu_ins.data_in[12] ),
    .B(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0530_));
 sky130_fd_sc_hd__nor2_1 _0957_ (.A(_0529_),
    .B(_0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0531_));
 sky130_fd_sc_hd__or4_1 _0958_ (.A(_0508_),
    .B(_0515_),
    .C(_0520_),
    .D(_0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0532_));
 sky130_fd_sc_hd__o41a_2 _0959_ (.A1(\dpu_ins.data_in[8] ),
    .A2(\dpu_ins.data_in[9] ),
    .A3(\dpu_ins.data_in[10] ),
    .A4(\dpu_ins.data_in[11] ),
    .B1(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0533_));
 sky130_fd_sc_hd__o21bai_1 _0960_ (.A1(_0505_),
    .A2(_0532_),
    .B1_N(_0533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0534_));
 sky130_fd_sc_hd__o21a_1 _0961_ (.A1(_0531_),
    .A2(_0534_),
    .B1(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0535_));
 sky130_fd_sc_hd__a21boi_1 _0962_ (.A1(_0531_),
    .A2(_0534_),
    .B1_N(_0535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0536_));
 sky130_fd_sc_hd__a221o_1 _0963_ (.A1(\dpu_ins.data_in[13] ),
    .A2(_0446_),
    .B1(_0462_),
    .B2(\dpu_ins.data_in[11] ),
    .C1(_0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[12] ));
 sky130_fd_sc_hd__a21oi_1 _0964_ (.A1(_0531_),
    .A2(_0534_),
    .B1(_0529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0537_));
 sky130_fd_sc_hd__and2_1 _0965_ (.A(\dpu_ins.data_in[13] ),
    .B(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0538_));
 sky130_fd_sc_hd__nor2_1 _0966_ (.A(\dpu_ins.data_in[13] ),
    .B(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0539_));
 sky130_fd_sc_hd__or2_1 _0967_ (.A(_0538_),
    .B(_0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0540_));
 sky130_fd_sc_hd__a21oi_1 _0968_ (.A1(_0537_),
    .A2(_0540_),
    .B1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0541_));
 sky130_fd_sc_hd__o21a_1 _0969_ (.A1(_0537_),
    .A2(_0540_),
    .B1(_0541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0542_));
 sky130_fd_sc_hd__a221o_1 _0970_ (.A1(\dpu_ins.data_in[14] ),
    .A2(_0446_),
    .B1(_0462_),
    .B2(\dpu_ins.data_in[12] ),
    .C1(_0542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[13] ));
 sky130_fd_sc_hd__nand2_1 _0971_ (.A(\dpu_ins.data_in[14] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0543_));
 sky130_fd_sc_hd__or2_1 _0972_ (.A(\dpu_ins.data_in[14] ),
    .B(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0544_));
 sky130_fd_sc_hd__nand2_1 _0973_ (.A(_0543_),
    .B(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0545_));
 sky130_fd_sc_hd__o21ba_1 _0974_ (.A1(_0537_),
    .A2(_0539_),
    .B1_N(_0538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0546_));
 sky130_fd_sc_hd__or2_1 _0975_ (.A(_0545_),
    .B(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0547_));
 sky130_fd_sc_hd__a21oi_1 _0976_ (.A1(_0545_),
    .A2(_0546_),
    .B1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0548_));
 sky130_fd_sc_hd__a22o_1 _0977_ (.A1(\dpu_ins.data_in[15] ),
    .A2(_0482_),
    .B1(_0483_),
    .B2(\dpu_ins.data_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0549_));
 sky130_fd_sc_hd__a21o_1 _0978_ (.A1(_0547_),
    .A2(_0548_),
    .B1(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[14] ));
 sky130_fd_sc_hd__buf_4 _0979_ (.A(_0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0550_));
 sky130_fd_sc_hd__buf_4 _0980_ (.A(_0461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0551_));
 sky130_fd_sc_hd__xnor2_1 _0981_ (.A(\dpu_ins.data_in[15] ),
    .B(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0552_));
 sky130_fd_sc_hd__a21oi_1 _0982_ (.A1(_0543_),
    .A2(_0547_),
    .B1(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0553_));
 sky130_fd_sc_hd__a31o_1 _0983_ (.A1(_0543_),
    .A2(_0547_),
    .A3(_0552_),
    .B1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0554_));
 sky130_fd_sc_hd__nor2_1 _0984_ (.A(_0553_),
    .B(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0555_));
 sky130_fd_sc_hd__a221o_1 _0985_ (.A1(\dpu_ins.data_in[16] ),
    .A2(_0550_),
    .B1(_0551_),
    .B2(\dpu_ins.data_in[14] ),
    .C1(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[15] ));
 sky130_fd_sc_hd__inv_2 _0986_ (.A(_0531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0556_));
 sky130_fd_sc_hd__or4_1 _0987_ (.A(_0556_),
    .B(_0540_),
    .C(_0545_),
    .D(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0557_));
 sky130_fd_sc_hd__nor3_1 _0988_ (.A(_0505_),
    .B(_0532_),
    .C(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0558_));
 sky130_fd_sc_hd__o41a_2 _0989_ (.A1(\dpu_ins.data_in[12] ),
    .A2(\dpu_ins.data_in[13] ),
    .A3(\dpu_ins.data_in[14] ),
    .A4(\dpu_ins.data_in[15] ),
    .B1(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0559_));
 sky130_fd_sc_hd__nor3_1 _0990_ (.A(_0533_),
    .B(net3),
    .C(_0559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2_1 _0991_ (.A(\dpu_ins.data_in[16] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0561_));
 sky130_fd_sc_hd__or2_1 _0992_ (.A(\dpu_ins.data_in[16] ),
    .B(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0562_));
 sky130_fd_sc_hd__nand2_1 _0993_ (.A(_0561_),
    .B(_0562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0563_));
 sky130_fd_sc_hd__nand2_1 _0994_ (.A(_0560_),
    .B(_0563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0564_));
 sky130_fd_sc_hd__or2_1 _0995_ (.A(_0560_),
    .B(_0563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0565_));
 sky130_fd_sc_hd__a22o_1 _0996_ (.A1(\dpu_ins.data_in[17] ),
    .A2(_0482_),
    .B1(_0483_),
    .B2(\dpu_ins.data_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0566_));
 sky130_fd_sc_hd__a31o_1 _0997_ (.A1(_0470_),
    .A2(_0564_),
    .A3(_0565_),
    .B1(_0566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[16] ));
 sky130_fd_sc_hd__xnor2_1 _0998_ (.A(\dpu_ins.data_in[17] ),
    .B(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0567_));
 sky130_fd_sc_hd__nand3_1 _0999_ (.A(_0561_),
    .B(_0565_),
    .C(_0567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0568_));
 sky130_fd_sc_hd__a21o_1 _1000_ (.A1(_0561_),
    .A2(_0565_),
    .B1(_0567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0569_));
 sky130_fd_sc_hd__a22o_1 _1001_ (.A1(\dpu_ins.data_in[18] ),
    .A2(_0482_),
    .B1(_0483_),
    .B2(\dpu_ins.data_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0570_));
 sky130_fd_sc_hd__a31o_1 _1002_ (.A1(_0470_),
    .A2(_0568_),
    .A3(_0569_),
    .B1(_0570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[17] ));
 sky130_fd_sc_hd__nand2_1 _1003_ (.A(\dpu_ins.data_in[18] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0571_));
 sky130_fd_sc_hd__or2_1 _1004_ (.A(\dpu_ins.data_in[18] ),
    .B(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0572_));
 sky130_fd_sc_hd__nand2_1 _1005_ (.A(_0571_),
    .B(_0572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0573_));
 sky130_fd_sc_hd__o21ai_1 _1006_ (.A1(\dpu_ins.data_in[16] ),
    .A2(\dpu_ins.data_in[17] ),
    .B1(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0574_));
 sky130_fd_sc_hd__a2bb2o_1 _1007_ (.A1_N(\dpu_ins.data_in[17] ),
    .A2_N(_0455_),
    .B1(_0565_),
    .B2(_0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0575_));
 sky130_fd_sc_hd__a21oi_1 _1008_ (.A1(_0573_),
    .A2(_0575_),
    .B1(\dpu_ins.cur_cmd[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0576_));
 sky130_fd_sc_hd__o21a_1 _1009_ (.A1(_0573_),
    .A2(_0575_),
    .B1(_0576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0577_));
 sky130_fd_sc_hd__a221o_1 _1010_ (.A1(\dpu_ins.data_in[19] ),
    .A2(_0550_),
    .B1(_0551_),
    .B2(\dpu_ins.data_in[17] ),
    .C1(_0577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[18] ));
 sky130_fd_sc_hd__nand2_1 _1011_ (.A(\dpu_ins.data_in[19] ),
    .B(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0578_));
 sky130_fd_sc_hd__or2_1 _1012_ (.A(\dpu_ins.data_in[19] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0579_));
 sky130_fd_sc_hd__nand2_1 _1013_ (.A(_0578_),
    .B(_0579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0580_));
 sky130_fd_sc_hd__o21ai_1 _1014_ (.A1(_0573_),
    .A2(_0575_),
    .B1(_0571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0581_));
 sky130_fd_sc_hd__xor2_1 _1015_ (.A(_0580_),
    .B(_0581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0582_));
 sky130_fd_sc_hd__nor2_1 _1016_ (.A(\dpu_ins.cur_cmd[6] ),
    .B(_0582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0583_));
 sky130_fd_sc_hd__a221o_1 _1017_ (.A1(\dpu_ins.data_in[20] ),
    .A2(_0550_),
    .B1(_0551_),
    .B2(\dpu_ins.data_in[18] ),
    .C1(_0583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[19] ));
 sky130_fd_sc_hd__nand3_1 _1018_ (.A(_0571_),
    .B(_0574_),
    .C(_0578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0584_));
 sky130_fd_sc_hd__or4_1 _1019_ (.A(_0563_),
    .B(_0567_),
    .C(_0573_),
    .D(_0580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0585_));
 sky130_fd_sc_hd__inv_2 _1020_ (.A(_0585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0586_));
 sky130_fd_sc_hd__o31a_1 _1021_ (.A1(_0533_),
    .A2(net3),
    .A3(_0559_),
    .B1(_0586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0587_));
 sky130_fd_sc_hd__and2_1 _1022_ (.A(\dpu_ins.data_in[20] ),
    .B(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0588_));
 sky130_fd_sc_hd__nor2_1 _1023_ (.A(\dpu_ins.data_in[20] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0589_));
 sky130_fd_sc_hd__or2_1 _1024_ (.A(_0588_),
    .B(_0589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0590_));
 sky130_fd_sc_hd__o21ba_1 _1025_ (.A1(_0584_),
    .A2(_0587_),
    .B1_N(_0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0591_));
 sky130_fd_sc_hd__or3b_1 _1026_ (.A(_0584_),
    .B(_0587_),
    .C_N(_0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0592_));
 sky130_fd_sc_hd__nor3b_1 _1027_ (.A(net12),
    .B(_0591_),
    .C_N(_0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0593_));
 sky130_fd_sc_hd__a221o_1 _1028_ (.A1(\dpu_ins.data_in[21] ),
    .A2(_0550_),
    .B1(_0551_),
    .B2(\dpu_ins.data_in[19] ),
    .C1(_0593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[20] ));
 sky130_fd_sc_hd__nor2_1 _1029_ (.A(_0588_),
    .B(_0591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0594_));
 sky130_fd_sc_hd__and2_1 _1030_ (.A(\dpu_ins.data_in[21] ),
    .B(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0595_));
 sky130_fd_sc_hd__nor2_1 _1031_ (.A(\dpu_ins.data_in[21] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0596_));
 sky130_fd_sc_hd__or2_1 _1032_ (.A(_0595_),
    .B(_0596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0597_));
 sky130_fd_sc_hd__a21oi_1 _1033_ (.A1(_0594_),
    .A2(_0597_),
    .B1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0598_));
 sky130_fd_sc_hd__o21a_1 _1034_ (.A1(_0594_),
    .A2(_0597_),
    .B1(_0598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0599_));
 sky130_fd_sc_hd__a221o_1 _1035_ (.A1(\dpu_ins.data_in[22] ),
    .A2(_0550_),
    .B1(_0551_),
    .B2(\dpu_ins.data_in[20] ),
    .C1(_0599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[21] ));
 sky130_fd_sc_hd__and2_1 _1036_ (.A(\dpu_ins.data_in[22] ),
    .B(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0600_));
 sky130_fd_sc_hd__nor2_1 _1037_ (.A(\dpu_ins.data_in[22] ),
    .B(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0601_));
 sky130_fd_sc_hd__nor2_1 _1038_ (.A(_0600_),
    .B(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_1 _1039_ (.A(\dpu_ins.data_in[21] ),
    .B(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0603_));
 sky130_fd_sc_hd__a21oi_1 _1040_ (.A1(_0603_),
    .A2(_0594_),
    .B1(_0596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0604_));
 sky130_fd_sc_hd__xnor2_1 _1041_ (.A(_0602_),
    .B(_0604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0605_));
 sky130_fd_sc_hd__nor2_1 _1042_ (.A(net12),
    .B(_0605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0606_));
 sky130_fd_sc_hd__a221o_1 _1043_ (.A1(\dpu_ins.data_in[23] ),
    .A2(_0550_),
    .B1(_0551_),
    .B2(\dpu_ins.data_in[21] ),
    .C1(_0606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[22] ));
 sky130_fd_sc_hd__xnor2_1 _1044_ (.A(\dpu_ins.data_in[23] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0607_));
 sky130_fd_sc_hd__a21oi_1 _1045_ (.A1(_0602_),
    .A2(_0604_),
    .B1(_0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0608_));
 sky130_fd_sc_hd__xor2_1 _1046_ (.A(_0607_),
    .B(_0608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0609_));
 sky130_fd_sc_hd__a22o_1 _1047_ (.A1(\dpu_ins.data_in[24] ),
    .A2(_0482_),
    .B1(_0483_),
    .B2(\dpu_ins.data_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0610_));
 sky130_fd_sc_hd__a21o_1 _1048_ (.A1(_0470_),
    .A2(_0609_),
    .B1(_0610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[23] ));
 sky130_fd_sc_hd__and3_1 _1049_ (.A(_0571_),
    .B(_0574_),
    .C(_0578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0611_));
 sky130_fd_sc_hd__a2111oi_1 _1050_ (.A1(\dpu_ins.data_in[23] ),
    .A2(_0454_),
    .B1(_0588_),
    .C1(_0595_),
    .D1(_0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0612_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(_0602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0613_));
 sky130_fd_sc_hd__nor4_1 _1052_ (.A(_0590_),
    .B(_0597_),
    .C(_0613_),
    .D(_0607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0614_));
 sky130_fd_sc_hd__o311ai_2 _1053_ (.A1(_0533_),
    .A2(net3),
    .A3(_0559_),
    .B1(_0586_),
    .C1(_0614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0615_));
 sky130_fd_sc_hd__nand3_1 _1054_ (.A(_0611_),
    .B(_0612_),
    .C(_0615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0616_));
 sky130_fd_sc_hd__nand2_1 _1055_ (.A(\dpu_ins.data_in[24] ),
    .B(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0617_));
 sky130_fd_sc_hd__or2_1 _1056_ (.A(\dpu_ins.data_in[24] ),
    .B(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0618_));
 sky130_fd_sc_hd__nand2_1 _1057_ (.A(_0617_),
    .B(_0618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0619_));
 sky130_fd_sc_hd__xnor2_1 _1058_ (.A(_0616_),
    .B(_0619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0620_));
 sky130_fd_sc_hd__a22o_1 _1059_ (.A1(\dpu_ins.data_in[25] ),
    .A2(_0482_),
    .B1(_0483_),
    .B2(\dpu_ins.data_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0621_));
 sky130_fd_sc_hd__a21o_1 _1060_ (.A1(_0470_),
    .A2(_0620_),
    .B1(_0621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[24] ));
 sky130_fd_sc_hd__a31o_1 _1061_ (.A1(_0611_),
    .A2(net4),
    .A3(_0615_),
    .B1(_0619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0622_));
 sky130_fd_sc_hd__and2_1 _1062_ (.A(\dpu_ins.data_in[25] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0623_));
 sky130_fd_sc_hd__nor2_1 _1063_ (.A(\dpu_ins.data_in[25] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0624_));
 sky130_fd_sc_hd__or2_1 _1064_ (.A(_0623_),
    .B(_0624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0625_));
 sky130_fd_sc_hd__a31o_1 _1065_ (.A1(_0617_),
    .A2(_0622_),
    .A3(_0625_),
    .B1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0626_));
 sky130_fd_sc_hd__a21o_1 _1066_ (.A1(_0617_),
    .A2(_0622_),
    .B1(_0625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0627_));
 sky130_fd_sc_hd__and2b_1 _1067_ (.A_N(_0626_),
    .B(_0627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0628_));
 sky130_fd_sc_hd__a221o_1 _1068_ (.A1(\dpu_ins.data_in[26] ),
    .A2(_0550_),
    .B1(_0551_),
    .B2(\dpu_ins.data_in[24] ),
    .C1(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[25] ));
 sky130_fd_sc_hd__nand2_1 _1069_ (.A(\dpu_ins.data_in[26] ),
    .B(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0629_));
 sky130_fd_sc_hd__or2_1 _1070_ (.A(\dpu_ins.data_in[26] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0630_));
 sky130_fd_sc_hd__nand2_1 _1071_ (.A(_0629_),
    .B(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0631_));
 sky130_fd_sc_hd__o21ai_1 _1072_ (.A1(\dpu_ins.data_in[24] ),
    .A2(\dpu_ins.data_in[25] ),
    .B1(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0632_));
 sky130_fd_sc_hd__a21o_1 _1073_ (.A1(_0622_),
    .A2(_0632_),
    .B1(_0624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0633_));
 sky130_fd_sc_hd__or2_1 _1074_ (.A(_0631_),
    .B(_0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0634_));
 sky130_fd_sc_hd__nand2_1 _1075_ (.A(_0631_),
    .B(_0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0635_));
 sky130_fd_sc_hd__a22o_1 _1076_ (.A1(\dpu_ins.data_in[27] ),
    .A2(_0482_),
    .B1(_0483_),
    .B2(\dpu_ins.data_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0636_));
 sky130_fd_sc_hd__a31o_1 _1077_ (.A1(_0470_),
    .A2(_0634_),
    .A3(_0635_),
    .B1(_0636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[26] ));
 sky130_fd_sc_hd__xnor2_1 _1078_ (.A(\dpu_ins.data_in[27] ),
    .B(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0637_));
 sky130_fd_sc_hd__a21oi_1 _1079_ (.A1(_0629_),
    .A2(_0634_),
    .B1(_0637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0638_));
 sky130_fd_sc_hd__a31o_1 _1080_ (.A1(_0629_),
    .A2(_0634_),
    .A3(_0637_),
    .B1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0639_));
 sky130_fd_sc_hd__nor2_1 _1081_ (.A(_0638_),
    .B(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0640_));
 sky130_fd_sc_hd__a221o_1 _1082_ (.A1(\dpu_ins.data_in[28] ),
    .A2(_0550_),
    .B1(_0551_),
    .B2(\dpu_ins.data_in[26] ),
    .C1(_0640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[27] ));
 sky130_fd_sc_hd__or3_1 _1083_ (.A(_0625_),
    .B(_0631_),
    .C(_0637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0641_));
 sky130_fd_sc_hd__o21ai_1 _1084_ (.A1(\dpu_ins.data_in[26] ),
    .A2(\dpu_ins.data_in[27] ),
    .B1(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0642_));
 sky130_fd_sc_hd__o211a_1 _1085_ (.A1(_0622_),
    .A2(_0641_),
    .B1(_0642_),
    .C1(_0632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0643_));
 sky130_fd_sc_hd__nand2_1 _1086_ (.A(\dpu_ins.data_in[28] ),
    .B(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0644_));
 sky130_fd_sc_hd__or2_1 _1087_ (.A(\dpu_ins.data_in[28] ),
    .B(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0645_));
 sky130_fd_sc_hd__nand2_1 _1088_ (.A(_0644_),
    .B(_0645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0646_));
 sky130_fd_sc_hd__a21oi_1 _1089_ (.A1(_0643_),
    .A2(_0646_),
    .B1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0647_));
 sky130_fd_sc_hd__o21a_1 _1090_ (.A1(_0643_),
    .A2(_0646_),
    .B1(_0647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0648_));
 sky130_fd_sc_hd__a221o_1 _1091_ (.A1(\dpu_ins.data_in[29] ),
    .A2(_0550_),
    .B1(_0551_),
    .B2(\dpu_ins.data_in[27] ),
    .C1(_0648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[28] ));
 sky130_fd_sc_hd__or2_1 _1092_ (.A(\dpu_ins.data_in[29] ),
    .B(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0649_));
 sky130_fd_sc_hd__nand2_1 _1093_ (.A(\dpu_ins.data_in[29] ),
    .B(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0650_));
 sky130_fd_sc_hd__nand2_1 _1094_ (.A(_0649_),
    .B(_0650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0651_));
 sky130_fd_sc_hd__o21a_1 _1095_ (.A1(_0643_),
    .A2(_0646_),
    .B1(_0644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0652_));
 sky130_fd_sc_hd__xnor2_1 _1096_ (.A(_0651_),
    .B(_0652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0653_));
 sky130_fd_sc_hd__nor2_1 _1097_ (.A(net12),
    .B(_0653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0654_));
 sky130_fd_sc_hd__a221o_1 _1098_ (.A1(\dpu_ins.data_in[30] ),
    .A2(_0550_),
    .B1(_0551_),
    .B2(\dpu_ins.data_in[28] ),
    .C1(_0654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[29] ));
 sky130_fd_sc_hd__or3_1 _1099_ (.A(_0643_),
    .B(_0646_),
    .C(_0651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0655_));
 sky130_fd_sc_hd__and2_1 _1100_ (.A(\dpu_ins.data_in[30] ),
    .B(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0656_));
 sky130_fd_sc_hd__nor2_1 _1101_ (.A(\dpu_ins.data_in[30] ),
    .B(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0657_));
 sky130_fd_sc_hd__or2_1 _1102_ (.A(_0656_),
    .B(_0657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0658_));
 sky130_fd_sc_hd__a31oi_2 _1103_ (.A1(_0644_),
    .A2(_0650_),
    .A3(_0655_),
    .B1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0659_));
 sky130_fd_sc_hd__a41o_1 _1104_ (.A1(_0644_),
    .A2(_0650_),
    .A3(_0658_),
    .A4(_0655_),
    .B1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0660_));
 sky130_fd_sc_hd__a22oi_1 _1105_ (.A1(\dpu_ins.data_in[31] ),
    .A2(_0482_),
    .B1(_0483_),
    .B2(\dpu_ins.data_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0661_));
 sky130_fd_sc_hd__o21ai_1 _1106_ (.A1(_0659_),
    .A2(_0660_),
    .B1(_0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(\dpu_ins.data_out[30] ));
 sky130_fd_sc_hd__xnor2_1 _1107_ (.A(\dpu_ins.data_in[31] ),
    .B(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0662_));
 sky130_fd_sc_hd__or3b_1 _1108_ (.A(_0656_),
    .B(_0659_),
    .C_N(_0662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0663_));
 sky130_fd_sc_hd__o21bai_1 _1109_ (.A1(_0656_),
    .A2(_0659_),
    .B1_N(_0662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0664_));
 sky130_fd_sc_hd__a32o_1 _1110_ (.A1(_0470_),
    .A2(_0663_),
    .A3(_0664_),
    .B1(net107),
    .B2(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.data_out[31] ));
 sky130_fd_sc_hd__inv_2 _1111_ (.A(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0665_));
 sky130_fd_sc_hd__or2b_2 _1112_ (.A(\SRAMController_ins.cur_state[2] ),
    .B_N(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0666_));
 sky130_fd_sc_hd__nand2_1 _1113_ (.A(net9),
    .B(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0667_));
 sky130_fd_sc_hd__o22a_1 _1114_ (.A1(_0417_),
    .A2(_0666_),
    .B1(_0667_),
    .B2(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0668_));
 sky130_fd_sc_hd__o21ai_1 _1115_ (.A1(net17),
    .A2(_0665_),
    .B1(_0668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0669_));
 sky130_fd_sc_hd__and3_1 _1116_ (.A(\SRAMController_ins.rx_valid ),
    .B(_0441_),
    .C(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0670_));
 sky130_fd_sc_hd__o21a_1 _1117_ (.A1(\SRAMController_ins.rx_data_out[7] ),
    .A2(\SRAMController_ins.rx_data_out[5] ),
    .B1(_0670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0671_));
 sky130_fd_sc_hd__clkbuf_4 _1118_ (.A(_0418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_4 _1119_ (.A(_0416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0673_));
 sky130_fd_sc_hd__or2_1 _1120_ (.A(_0413_),
    .B(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _1121_ (.A0(_0672_),
    .A1(_0674_),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0675_));
 sky130_fd_sc_hd__and2b_1 _1122_ (.A_N(\SRAMController_ins.cur_state[0] ),
    .B(\SRAMController_ins.cur_state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_1 _1123_ (.A(net7),
    .B(_0676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0677_));
 sky130_fd_sc_hd__and2b_1 _1124_ (.A_N(\SRAMController_ins.cur_state[2] ),
    .B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0678_));
 sky130_fd_sc_hd__and3b_1 _1125_ (.A_N(net8),
    .B(\SRAMController_ins.cur_state[0] ),
    .C(_0678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0679_));
 sky130_fd_sc_hd__a22o_1 _1126_ (.A1(net8),
    .A2(_0415_),
    .B1(_0442_),
    .B2(_0678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _1127_ (.A0(_0679_),
    .A1(_0680_),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0681_));
 sky130_fd_sc_hd__o21bai_1 _1128_ (.A1(net8),
    .A2(_0677_),
    .B1_N(_0681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0682_));
 sky130_fd_sc_hd__or4_1 _1129_ (.A(_0669_),
    .B(_0671_),
    .C(_0675_),
    .D(_0682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_1 _1130_ (.A(_0683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.nxt_state[0] ));
 sky130_fd_sc_hd__inv_2 _1131_ (.A(\SRAMController_ins.rx_data_out[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_2 _1132_ (.A(net18),
    .B(\SRAMController_ins.uart_ready ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0685_));
 sky130_fd_sc_hd__a21oi_1 _1133_ (.A1(_0684_),
    .A2(\SRAMController_ins.rx_data_out[5] ),
    .B1(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0686_));
 sky130_fd_sc_hd__nor2_1 _1134_ (.A(net8),
    .B(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0687_));
 sky130_fd_sc_hd__or2_1 _1135_ (.A(_0411_),
    .B(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0688_));
 sky130_fd_sc_hd__and3_1 _1136_ (.A(net17),
    .B(net9),
    .C(\SRAMController_ins.cur_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0689_));
 sky130_fd_sc_hd__a2bb2o_1 _1137_ (.A1_N(_0688_),
    .A2_N(_0689_),
    .B1(net18),
    .B2(_0679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0690_));
 sky130_fd_sc_hd__a221o_1 _1138_ (.A1(net8),
    .A2(_0415_),
    .B1(_0687_),
    .B2(net7),
    .C1(_0690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0691_));
 sky130_fd_sc_hd__or3b_1 _1139_ (.A(_0686_),
    .B(_0691_),
    .C_N(_0668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_1 _1140_ (.A(_0692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.nxt_state[1] ));
 sky130_fd_sc_hd__nor3_1 _1141_ (.A(\SRAMController_ins.rx_data_out[7] ),
    .B(\SRAMController_ins.rx_data_out[5] ),
    .C(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0693_));
 sky130_fd_sc_hd__and3_1 _1142_ (.A(\SRAMController_ins.cur_state[2] ),
    .B(\SRAMController_ins.cur_state[3] ),
    .C(_0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0694_));
 sky130_fd_sc_hd__a2111o_1 _1143_ (.A1(net17),
    .A2(_0672_),
    .B1(_0693_),
    .C1(_0694_),
    .D1(_0415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0695_));
 sky130_fd_sc_hd__or2_1 _1144_ (.A(_0669_),
    .B(_0695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0696_));
 sky130_fd_sc_hd__clkbuf_1 _1145_ (.A(_0696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.nxt_state[2] ));
 sky130_fd_sc_hd__inv_2 _1146_ (.A(_0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0697_));
 sky130_fd_sc_hd__nor2_4 _1147_ (.A(_0684_),
    .B(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0698_));
 sky130_fd_sc_hd__a221o_1 _1148_ (.A1(\SRAMController_ins.cur_state[3] ),
    .A2(_0412_),
    .B1(_0697_),
    .B2(net18),
    .C1(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.nxt_state[3] ));
 sky130_fd_sc_hd__nor2_8 _1149_ (.A(_0412_),
    .B(_0666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0699_));
 sky130_fd_sc_hd__and3_1 _1150_ (.A(net8),
    .B(net7),
    .C(_0676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0700_));
 sky130_fd_sc_hd__buf_4 _1151_ (.A(_0700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0701_));
 sky130_fd_sc_hd__a31o_1 _1152_ (.A1(net9),
    .A2(\SRAMController_ins.cur_state[0] ),
    .A3(_0678_),
    .B1(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0702_));
 sky130_fd_sc_hd__and3_1 _1153_ (.A(_0684_),
    .B(\SRAMController_ins.rx_data_out[5] ),
    .C(_0670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0703_));
 sky130_fd_sc_hd__and2_1 _1154_ (.A(\SRAMController_ins.rx_data_out[0] ),
    .B(_0703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0704_));
 sky130_fd_sc_hd__a221o_1 _1155_ (.A1(\SRAMController_ins.addr_tmp[0] ),
    .A2(_0699_),
    .B1(_0702_),
    .B2(\SRAMController_ins.sram_addr_from_dpu[0] ),
    .C1(_0704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.addr[0] ));
 sky130_fd_sc_hd__and2_1 _1156_ (.A(\SRAMController_ins.rx_data_out[1] ),
    .B(_0703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0705_));
 sky130_fd_sc_hd__a221o_1 _1157_ (.A1(\SRAMController_ins.addr_tmp[1] ),
    .A2(_0699_),
    .B1(_0702_),
    .B2(\SRAMController_ins.sram_addr_from_dpu[1] ),
    .C1(_0705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.addr[1] ));
 sky130_fd_sc_hd__and2_1 _1158_ (.A(\SRAMController_ins.rx_data_out[2] ),
    .B(_0703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0706_));
 sky130_fd_sc_hd__a221o_1 _1159_ (.A1(\SRAMController_ins.addr_tmp[2] ),
    .A2(_0699_),
    .B1(_0702_),
    .B2(\SRAMController_ins.sram_addr_from_dpu[2] ),
    .C1(_0706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.addr[2] ));
 sky130_fd_sc_hd__and2_1 _1160_ (.A(\SRAMController_ins.rx_data_out[3] ),
    .B(_0703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0707_));
 sky130_fd_sc_hd__a221o_1 _1161_ (.A1(\SRAMController_ins.addr_tmp[3] ),
    .A2(_0699_),
    .B1(_0702_),
    .B2(\SRAMController_ins.sram_addr_from_dpu[3] ),
    .C1(_0707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.addr[3] ));
 sky130_fd_sc_hd__a31o_1 _1162_ (.A1(net8),
    .A2(\SRAMController_ins.cur_state[0] ),
    .A3(_0678_),
    .B1(_0703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.we_n ));
 sky130_fd_sc_hd__a31o_1 _1163_ (.A1(_0684_),
    .A2(\SRAMController_ins.rx_data_out[5] ),
    .A3(net18),
    .B1(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0708_));
 sky130_fd_sc_hd__or4b_1 _1164_ (.A(_0420_),
    .B(_0679_),
    .C(_0694_),
    .D_N(_0708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0709_));
 sky130_fd_sc_hd__or2b_1 _1165_ (.A(_0673_),
    .B_N(_0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0710_));
 sky130_fd_sc_hd__or3_1 _1166_ (.A(_0680_),
    .B(_0709_),
    .C(_0710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0711_));
 sky130_fd_sc_hd__buf_1 _1167_ (.A(_0711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.csb_n ));
 sky130_fd_sc_hd__mux2_1 _1168_ (.A0(\dpu_ins.cur_state[1] ),
    .A1(_0677_),
    .S(\dpu_ins.cur_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0712_));
 sky130_fd_sc_hd__or2_1 _1169_ (.A(_0698_),
    .B(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0713_));
 sky130_fd_sc_hd__clkbuf_1 _1170_ (.A(_0713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\dpu_ins.nxt_state[0] ));
 sky130_fd_sc_hd__or3b_1 _1171_ (.A(\dpu_ins.cur_state[1] ),
    .B(_0677_),
    .C_N(\dpu_ins.cur_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0714_));
 sky130_fd_sc_hd__buf_4 _1172_ (.A(_0714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0715_));
 sky130_fd_sc_hd__clkbuf_4 _1173_ (.A(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0716_));
 sky130_fd_sc_hd__and2_1 _1174_ (.A(net7),
    .B(_0676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0717_));
 sky130_fd_sc_hd__a21bo_1 _1175_ (.A1(\dpu_ins.cur_state[0] ),
    .A2(_0717_),
    .B1_N(\dpu_ins.cur_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0718_));
 sky130_fd_sc_hd__nand2_1 _1176_ (.A(_0716_),
    .B(_0718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(\dpu_ins.nxt_state[1] ));
 sky130_fd_sc_hd__buf_2 _1177_ (.A(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0719_));
 sky130_fd_sc_hd__buf_2 _1178_ (.A(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0720_));
 sky130_fd_sc_hd__a22o_1 _1179_ (.A1(\SRAMController_ins.data_tmp[0] ),
    .A2(_0719_),
    .B1(_0720_),
    .B2(\SRAMController_ins.sram_data_from_dpu[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[0] ));
 sky130_fd_sc_hd__a22o_1 _1180_ (.A1(\SRAMController_ins.data_tmp[1] ),
    .A2(_0719_),
    .B1(_0720_),
    .B2(\SRAMController_ins.sram_data_from_dpu[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[1] ));
 sky130_fd_sc_hd__a22o_1 _1181_ (.A1(\SRAMController_ins.data_tmp[2] ),
    .A2(_0719_),
    .B1(_0720_),
    .B2(\SRAMController_ins.sram_data_from_dpu[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[2] ));
 sky130_fd_sc_hd__a22o_1 _1182_ (.A1(\SRAMController_ins.data_tmp[3] ),
    .A2(_0719_),
    .B1(_0720_),
    .B2(\SRAMController_ins.sram_data_from_dpu[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[3] ));
 sky130_fd_sc_hd__a22o_1 _1183_ (.A1(\SRAMController_ins.data_tmp[4] ),
    .A2(_0719_),
    .B1(_0720_),
    .B2(\SRAMController_ins.sram_data_from_dpu[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[4] ));
 sky130_fd_sc_hd__a22o_1 _1184_ (.A1(\SRAMController_ins.data_tmp[5] ),
    .A2(_0719_),
    .B1(_0720_),
    .B2(\SRAMController_ins.sram_data_from_dpu[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[5] ));
 sky130_fd_sc_hd__a22o_1 _1185_ (.A1(\SRAMController_ins.data_tmp[6] ),
    .A2(_0719_),
    .B1(_0720_),
    .B2(\SRAMController_ins.sram_data_from_dpu[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[6] ));
 sky130_fd_sc_hd__a22o_1 _1186_ (.A1(\SRAMController_ins.data_tmp[7] ),
    .A2(_0719_),
    .B1(_0720_),
    .B2(\SRAMController_ins.sram_data_from_dpu[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[7] ));
 sky130_fd_sc_hd__a22o_1 _1187_ (.A1(\SRAMController_ins.data_tmp[8] ),
    .A2(_0719_),
    .B1(_0720_),
    .B2(\SRAMController_ins.sram_data_from_dpu[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[8] ));
 sky130_fd_sc_hd__a22o_1 _1188_ (.A1(\SRAMController_ins.data_tmp[9] ),
    .A2(_0719_),
    .B1(_0720_),
    .B2(\SRAMController_ins.sram_data_from_dpu[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[9] ));
 sky130_fd_sc_hd__buf_2 _1189_ (.A(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0721_));
 sky130_fd_sc_hd__buf_2 _1190_ (.A(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0722_));
 sky130_fd_sc_hd__a22o_1 _1191_ (.A1(\SRAMController_ins.data_tmp[10] ),
    .A2(_0721_),
    .B1(_0722_),
    .B2(\SRAMController_ins.sram_data_from_dpu[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[10] ));
 sky130_fd_sc_hd__a22o_1 _1192_ (.A1(\SRAMController_ins.data_tmp[11] ),
    .A2(_0721_),
    .B1(_0722_),
    .B2(\SRAMController_ins.sram_data_from_dpu[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[11] ));
 sky130_fd_sc_hd__a22o_1 _1193_ (.A1(\SRAMController_ins.data_tmp[12] ),
    .A2(_0721_),
    .B1(_0722_),
    .B2(\SRAMController_ins.sram_data_from_dpu[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[12] ));
 sky130_fd_sc_hd__a22o_1 _1194_ (.A1(\SRAMController_ins.data_tmp[13] ),
    .A2(_0721_),
    .B1(_0722_),
    .B2(\SRAMController_ins.sram_data_from_dpu[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[13] ));
 sky130_fd_sc_hd__a22o_1 _1195_ (.A1(\SRAMController_ins.data_tmp[14] ),
    .A2(_0721_),
    .B1(_0722_),
    .B2(\SRAMController_ins.sram_data_from_dpu[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[14] ));
 sky130_fd_sc_hd__a22o_1 _1196_ (.A1(\SRAMController_ins.data_tmp[15] ),
    .A2(_0721_),
    .B1(_0722_),
    .B2(\SRAMController_ins.sram_data_from_dpu[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[15] ));
 sky130_fd_sc_hd__a22o_1 _1197_ (.A1(\SRAMController_ins.data_tmp[16] ),
    .A2(_0721_),
    .B1(_0722_),
    .B2(\SRAMController_ins.sram_data_from_dpu[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[16] ));
 sky130_fd_sc_hd__a22o_1 _1198_ (.A1(\SRAMController_ins.data_tmp[17] ),
    .A2(_0721_),
    .B1(_0722_),
    .B2(\SRAMController_ins.sram_data_from_dpu[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[17] ));
 sky130_fd_sc_hd__a22o_1 _1199_ (.A1(\SRAMController_ins.data_tmp[18] ),
    .A2(_0721_),
    .B1(_0722_),
    .B2(\SRAMController_ins.sram_data_from_dpu[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[18] ));
 sky130_fd_sc_hd__a22o_1 _1200_ (.A1(\SRAMController_ins.data_tmp[19] ),
    .A2(_0721_),
    .B1(_0722_),
    .B2(\SRAMController_ins.sram_data_from_dpu[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[19] ));
 sky130_fd_sc_hd__buf_2 _1201_ (.A(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0723_));
 sky130_fd_sc_hd__buf_2 _1202_ (.A(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0724_));
 sky130_fd_sc_hd__a22o_1 _1203_ (.A1(\SRAMController_ins.data_tmp[20] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(\SRAMController_ins.sram_data_from_dpu[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[20] ));
 sky130_fd_sc_hd__a22o_1 _1204_ (.A1(\SRAMController_ins.data_tmp[21] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(\SRAMController_ins.sram_data_from_dpu[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[21] ));
 sky130_fd_sc_hd__a22o_1 _1205_ (.A1(\SRAMController_ins.data_tmp[22] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(\SRAMController_ins.sram_data_from_dpu[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[22] ));
 sky130_fd_sc_hd__a22o_1 _1206_ (.A1(\SRAMController_ins.data_tmp[23] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(\SRAMController_ins.sram_data_from_dpu[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[23] ));
 sky130_fd_sc_hd__a22o_1 _1207_ (.A1(\SRAMController_ins.data_tmp[24] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(\SRAMController_ins.sram_data_from_dpu[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[24] ));
 sky130_fd_sc_hd__a22o_1 _1208_ (.A1(\SRAMController_ins.data_tmp[25] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(\SRAMController_ins.sram_data_from_dpu[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[25] ));
 sky130_fd_sc_hd__a22o_1 _1209_ (.A1(\SRAMController_ins.data_tmp[26] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(\SRAMController_ins.sram_data_from_dpu[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[26] ));
 sky130_fd_sc_hd__a22o_1 _1210_ (.A1(\SRAMController_ins.data_tmp[27] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(\SRAMController_ins.sram_data_from_dpu[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[27] ));
 sky130_fd_sc_hd__a22o_1 _1211_ (.A1(\SRAMController_ins.data_tmp[28] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(\SRAMController_ins.sram_data_from_dpu[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[28] ));
 sky130_fd_sc_hd__a22o_1 _1212_ (.A1(\SRAMController_ins.data_tmp[29] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(\SRAMController_ins.sram_data_from_dpu[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[29] ));
 sky130_fd_sc_hd__a22o_1 _1213_ (.A1(\SRAMController_ins.data_tmp[30] ),
    .A2(_0699_),
    .B1(_0701_),
    .B2(\SRAMController_ins.sram_data_from_dpu[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[30] ));
 sky130_fd_sc_hd__a22o_1 _1214_ (.A1(\SRAMController_ins.data_tmp[31] ),
    .A2(_0699_),
    .B1(_0701_),
    .B2(\SRAMController_ins.sram_data_from_dpu[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[31] ));
 sky130_fd_sc_hd__nand2_1 _1215_ (.A(net18),
    .B(_0437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0725_));
 sky130_fd_sc_hd__inv_2 _1216_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0726_));
 sky130_fd_sc_hd__a21oi_1 _1217_ (.A1(_0726_),
    .A2(_0403_),
    .B1(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0727_));
 sky130_fd_sc_hd__o21ai_1 _1218_ (.A1(_0437_),
    .A2(_0727_),
    .B1(_0435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0728_));
 sky130_fd_sc_hd__inv_2 _1219_ (.A(_0728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0729_));
 sky130_fd_sc_hd__nand2_1 _1220_ (.A(_0725_),
    .B(_0729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0730_));
 sky130_fd_sc_hd__mux2_1 _1221_ (.A0(net14),
    .A1(\UARTReceiver_ins.out_latched ),
    .S(_0730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0731_));
 sky130_fd_sc_hd__and3_1 _1222_ (.A(net28),
    .B(_0384_),
    .C(_0731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0732_));
 sky130_fd_sc_hd__clkbuf_1 _1223_ (.A(_0732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0008_));
 sky130_fd_sc_hd__o211a_1 _1224_ (.A1(_0399_),
    .A2(_0387_),
    .B1(_0435_),
    .C1(_0384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0733_));
 sky130_fd_sc_hd__nand2b_4 _1225_ (.A_N(net14),
    .B(_0733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0734_));
 sky130_fd_sc_hd__o31a_1 _1226_ (.A1(\UARTReceiver_ins.bitIndex[2] ),
    .A2(\UARTReceiver_ins.bitIndex[1] ),
    .A3(\UARTReceiver_ins.bitIndex[0] ),
    .B1(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0735_));
 sky130_fd_sc_hd__o21ai_1 _1227_ (.A1(_0734_),
    .A2(_0735_),
    .B1(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0736_));
 sky130_fd_sc_hd__nor2_1 _1228_ (.A(\UARTReceiver_ins.inputReg[1] ),
    .B(\UARTReceiver_ins.inputReg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0737_));
 sky130_fd_sc_hd__nor2_1 _1229_ (.A(\UARTReceiver_ins.inputReg[2] ),
    .B(_0385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0738_));
 sky130_fd_sc_hd__or4_4 _1230_ (.A(_0399_),
    .B(_0737_),
    .C(_0734_),
    .D(_0738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0739_));
 sky130_fd_sc_hd__or4_1 _1231_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .B(net19),
    .C(\UARTReceiver_ins.bitIndex[0] ),
    .D(_0739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0740_));
 sky130_fd_sc_hd__a21oi_1 _1232_ (.A1(_0736_),
    .A2(_0740_),
    .B1(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0009_));
 sky130_fd_sc_hd__or3b_1 _1233_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .B(net19),
    .C_N(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0741_));
 sky130_fd_sc_hd__and2_1 _1234_ (.A(net15),
    .B(_0741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0742_));
 sky130_fd_sc_hd__o21a_1 _1235_ (.A1(_0734_),
    .A2(_0742_),
    .B1(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0743_));
 sky130_fd_sc_hd__nor2_1 _1236_ (.A(_0739_),
    .B(_0741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0744_));
 sky130_fd_sc_hd__o21a_1 _1237_ (.A1(_0743_),
    .A2(_0744_),
    .B1(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0010_));
 sky130_fd_sc_hd__inv_2 _1238_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0745_));
 sky130_fd_sc_hd__and2b_1 _1239_ (.A_N(net20),
    .B(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0746_));
 sky130_fd_sc_hd__nand2_1 _1240_ (.A(_0745_),
    .B(_0746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0747_));
 sky130_fd_sc_hd__and2_1 _1241_ (.A(net15),
    .B(_0747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0748_));
 sky130_fd_sc_hd__o21a_1 _1242_ (.A1(_0734_),
    .A2(_0748_),
    .B1(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0749_));
 sky130_fd_sc_hd__nor2_1 _1243_ (.A(_0739_),
    .B(_0747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0750_));
 sky130_fd_sc_hd__o21a_1 _1244_ (.A1(_0749_),
    .A2(_0750_),
    .B1(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0011_));
 sky130_fd_sc_hd__inv_2 _1245_ (.A(_0739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0751_));
 sky130_fd_sc_hd__a31oi_1 _1246_ (.A1(_0745_),
    .A2(net19),
    .A3(net20),
    .B1(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0752_));
 sky130_fd_sc_hd__o21a_1 _1247_ (.A1(_0734_),
    .A2(_0752_),
    .B1(\UARTReceiver_ins.data[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0753_));
 sky130_fd_sc_hd__a41o_1 _1248_ (.A1(_0745_),
    .A2(net19),
    .A3(net20),
    .A4(_0751_),
    .B1(_0753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0754_));
 sky130_fd_sc_hd__and2_1 _1249_ (.A(net22),
    .B(_0754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0755_));
 sky130_fd_sc_hd__clkbuf_1 _1250_ (.A(_0755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0012_));
 sky130_fd_sc_hd__or3_1 _1251_ (.A(_0745_),
    .B(net19),
    .C(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0756_));
 sky130_fd_sc_hd__and2_1 _1252_ (.A(net15),
    .B(_0756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0757_));
 sky130_fd_sc_hd__o21a_1 _1253_ (.A1(_0734_),
    .A2(_0757_),
    .B1(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0758_));
 sky130_fd_sc_hd__nor2_1 _1254_ (.A(_0739_),
    .B(_0756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0759_));
 sky130_fd_sc_hd__o21a_1 _1255_ (.A1(_0758_),
    .A2(_0759_),
    .B1(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0013_));
 sky130_fd_sc_hd__and2b_1 _1256_ (.A_N(net19),
    .B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0760_));
 sky130_fd_sc_hd__a21oi_1 _1257_ (.A1(\UARTReceiver_ins.bitIndex[2] ),
    .A2(_0760_),
    .B1(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0761_));
 sky130_fd_sc_hd__o21a_1 _1258_ (.A1(_0734_),
    .A2(_0761_),
    .B1(\UARTReceiver_ins.data[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0762_));
 sky130_fd_sc_hd__a31o_1 _1259_ (.A1(\UARTReceiver_ins.bitIndex[2] ),
    .A2(_0751_),
    .A3(_0760_),
    .B1(_0762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0763_));
 sky130_fd_sc_hd__and2_1 _1260_ (.A(net22),
    .B(_0763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0764_));
 sky130_fd_sc_hd__clkbuf_1 _1261_ (.A(_0764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0014_));
 sky130_fd_sc_hd__a21oi_1 _1262_ (.A1(\UARTReceiver_ins.bitIndex[2] ),
    .A2(_0746_),
    .B1(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0765_));
 sky130_fd_sc_hd__o21a_1 _1263_ (.A1(_0734_),
    .A2(_0765_),
    .B1(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0766_));
 sky130_fd_sc_hd__and3_1 _1264_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .B(_0751_),
    .C(_0746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0767_));
 sky130_fd_sc_hd__o21a_1 _1265_ (.A1(_0766_),
    .A2(_0767_),
    .B1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0015_));
 sky130_fd_sc_hd__a21o_1 _1266_ (.A1(\UARTReceiver_ins.state[1] ),
    .A2(_0400_),
    .B1(_0734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0768_));
 sky130_fd_sc_hd__o2bb2a_1 _1267_ (.A1_N(\UARTReceiver_ins.data[7] ),
    .A2_N(_0768_),
    .B1(_0739_),
    .B2(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0769_));
 sky130_fd_sc_hd__nor2_1 _1268_ (.A(_0398_),
    .B(_0769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0016_));
 sky130_fd_sc_hd__nor2_2 _1269_ (.A(net14),
    .B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0770_));
 sky130_fd_sc_hd__a311oi_4 _1270_ (.A1(_0726_),
    .A2(_0403_),
    .A3(_0770_),
    .B1(net6),
    .C1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0771_));
 sky130_fd_sc_hd__and2_1 _1271_ (.A(\UARTReceiver_ins.sampleCount[0] ),
    .B(_0771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0772_));
 sky130_fd_sc_hd__a31oi_2 _1272_ (.A1(_0435_),
    .A2(_0770_),
    .A3(_0771_),
    .B1(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0773_));
 sky130_fd_sc_hd__or2_1 _1273_ (.A(\UARTReceiver_ins.sampleCount[0] ),
    .B(_0771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0774_));
 sky130_fd_sc_hd__and3b_1 _1274_ (.A_N(_0772_),
    .B(_0773_),
    .C(_0774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0775_));
 sky130_fd_sc_hd__clkbuf_1 _1275_ (.A(_0775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0017_));
 sky130_fd_sc_hd__nand2_1 _1276_ (.A(\UARTReceiver_ins.sampleCount[1] ),
    .B(_0772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0776_));
 sky130_fd_sc_hd__o211a_1 _1277_ (.A1(\UARTReceiver_ins.sampleCount[1] ),
    .A2(_0772_),
    .B1(_0776_),
    .C1(_0773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0018_));
 sky130_fd_sc_hd__a31o_1 _1278_ (.A1(\UARTReceiver_ins.sampleCount[1] ),
    .A2(\UARTReceiver_ins.sampleCount[0] ),
    .A3(_0771_),
    .B1(\UARTReceiver_ins.sampleCount[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0777_));
 sky130_fd_sc_hd__nand3_1 _1279_ (.A(\UARTReceiver_ins.sampleCount[2] ),
    .B(\UARTReceiver_ins.sampleCount[1] ),
    .C(_0772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0778_));
 sky130_fd_sc_hd__and3_1 _1280_ (.A(_0773_),
    .B(_0777_),
    .C(_0778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0779_));
 sky130_fd_sc_hd__clkbuf_1 _1281_ (.A(_0779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0019_));
 sky130_fd_sc_hd__inv_2 _1282_ (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0780_));
 sky130_fd_sc_hd__o21a_1 _1283_ (.A1(_0387_),
    .A2(_0770_),
    .B1(_0771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0177_));
 sky130_fd_sc_hd__a211oi_1 _1284_ (.A1(_0780_),
    .A2(_0778_),
    .B1(_0177_),
    .C1(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0020_));
 sky130_fd_sc_hd__o32a_1 _1285_ (.A1(net16),
    .A2(net2),
    .A3(_0390_),
    .B1(_0389_),
    .B2(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0021_));
 sky130_fd_sc_hd__o32a_1 _1286_ (.A1(net90),
    .A2(net16),
    .A3(_0390_),
    .B1(_0389_),
    .B2(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0022_));
 sky130_fd_sc_hd__o32a_1 _1287_ (.A1(net117),
    .A2(net16),
    .A3(_0390_),
    .B1(_0389_),
    .B2(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _1288_ (.A(net15),
    .B(_0733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0178_));
 sky130_fd_sc_hd__o31a_1 _1289_ (.A1(net16),
    .A2(\UARTReceiver_ins.state[2] ),
    .A3(net15),
    .B1(_0733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_1 _1290_ (.A(net20),
    .B(_0179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0180_));
 sky130_fd_sc_hd__o211a_1 _1291_ (.A1(net20),
    .A2(_0178_),
    .B1(_0180_),
    .C1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0024_));
 sky130_fd_sc_hd__o31ai_1 _1292_ (.A1(net16),
    .A2(\UARTReceiver_ins.state[2] ),
    .A3(net15),
    .B1(_0733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0181_));
 sky130_fd_sc_hd__or2_1 _1293_ (.A(_0760_),
    .B(_0746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0182_));
 sky130_fd_sc_hd__a22o_1 _1294_ (.A1(net19),
    .A2(_0181_),
    .B1(_0182_),
    .B2(_0178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0183_));
 sky130_fd_sc_hd__and2_1 _1295_ (.A(net25),
    .B(_0183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _1296_ (.A(_0184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0025_));
 sky130_fd_sc_hd__a31o_1 _1297_ (.A1(net19),
    .A2(net20),
    .A3(_0179_),
    .B1(\UARTReceiver_ins.bitIndex[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0185_));
 sky130_fd_sc_hd__a21o_1 _1298_ (.A1(net15),
    .A2(_0400_),
    .B1(_0181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _1299_ (.A(net25),
    .B(_0185_),
    .C(_0186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_1 _1300_ (.A(_0187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _1301_ (.A0(\SRAMController_ins.addr_tmp[0] ),
    .A1(\SRAMController_ins.rx_data_out[0] ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _1302_ (.A(_0188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1303_ (.A0(\SRAMController_ins.addr_tmp[1] ),
    .A1(\SRAMController_ins.rx_data_out[1] ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_1 _1304_ (.A(_0189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1305_ (.A0(\SRAMController_ins.addr_tmp[2] ),
    .A1(\SRAMController_ins.rx_data_out[2] ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_1 _1306_ (.A(_0190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1307_ (.A0(\SRAMController_ins.addr_tmp[3] ),
    .A1(\SRAMController_ins.rx_data_out[3] ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_1 _1308_ (.A(_0191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0030_));
 sky130_fd_sc_hd__a31o_1 _1309_ (.A1(net18),
    .A2(_0384_),
    .A3(_0729_),
    .B1(\UARTReceiver_ins.overrun ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0192_));
 sky130_fd_sc_hd__or3_1 _1310_ (.A(net14),
    .B(_0388_),
    .C(_0728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0193_));
 sky130_fd_sc_hd__and3_1 _1311_ (.A(net28),
    .B(_0192_),
    .C(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _1312_ (.A(_0194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0031_));
 sky130_fd_sc_hd__a21oi_1 _1313_ (.A1(net13),
    .A2(_0387_),
    .B1(_0727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _1314_ (.A(\UARTReceiver_ins.error ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0196_));
 sky130_fd_sc_hd__o41ai_1 _1315_ (.A1(_0388_),
    .A2(_0436_),
    .A3(_0439_),
    .A4(_0195_),
    .B1(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0197_));
 sky130_fd_sc_hd__and3_1 _1316_ (.A(net28),
    .B(_0193_),
    .C(_0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _1317_ (.A(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0032_));
 sky130_fd_sc_hd__o21a_1 _1318_ (.A1(net16),
    .A2(_0388_),
    .B1(\UARTReceiver_ins.out_latched ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0199_));
 sky130_fd_sc_hd__a31o_1 _1319_ (.A1(net8),
    .A2(net7),
    .A3(_0414_),
    .B1(_0710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0200_));
 sky130_fd_sc_hd__o41a_1 _1320_ (.A1(\UARTReceiver_ins.out_latched ),
    .A2(_0687_),
    .A3(_0717_),
    .A4(_0200_),
    .B1(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0201_));
 sky130_fd_sc_hd__nor2_1 _1321_ (.A(net16),
    .B(_0390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0202_));
 sky130_fd_sc_hd__o22a_1 _1322_ (.A1(net18),
    .A2(_0199_),
    .B1(_0201_),
    .B2(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0033_));
 sky130_fd_sc_hd__and2b_1 _1323_ (.A_N(net13),
    .B(\UARTReceiver_ins.state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0203_));
 sky130_fd_sc_hd__o211a_2 _1324_ (.A1(_0437_),
    .A2(_0203_),
    .B1(_0725_),
    .C1(_0384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0204_));
 sky130_fd_sc_hd__nor2_2 _1325_ (.A(_0398_),
    .B(_0204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0205_));
 sky130_fd_sc_hd__and3_1 _1326_ (.A(net13),
    .B(\UARTReceiver_ins.data[0] ),
    .C(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0206_));
 sky130_fd_sc_hd__o22a_1 _1327_ (.A1(\SRAMController_ins.rx_data_out[0] ),
    .A2(_0204_),
    .B1(_0205_),
    .B2(_0206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0034_));
 sky130_fd_sc_hd__and3_1 _1328_ (.A(net13),
    .B(\UARTReceiver_ins.data[1] ),
    .C(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0207_));
 sky130_fd_sc_hd__o22a_1 _1329_ (.A1(\SRAMController_ins.rx_data_out[1] ),
    .A2(_0204_),
    .B1(_0205_),
    .B2(_0207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0035_));
 sky130_fd_sc_hd__and3_1 _1330_ (.A(net13),
    .B(\UARTReceiver_ins.data[2] ),
    .C(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0208_));
 sky130_fd_sc_hd__o22a_1 _1331_ (.A1(\SRAMController_ins.rx_data_out[2] ),
    .A2(_0204_),
    .B1(_0205_),
    .B2(_0208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0036_));
 sky130_fd_sc_hd__and3_1 _1332_ (.A(net13),
    .B(\UARTReceiver_ins.data[3] ),
    .C(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0209_));
 sky130_fd_sc_hd__o22a_1 _1333_ (.A1(\SRAMController_ins.rx_data_out[3] ),
    .A2(_0204_),
    .B1(_0205_),
    .B2(_0209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0037_));
 sky130_fd_sc_hd__and3_1 _1334_ (.A(net13),
    .B(\UARTReceiver_ins.data[4] ),
    .C(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0210_));
 sky130_fd_sc_hd__o22a_1 _1335_ (.A1(net99),
    .A2(_0204_),
    .B1(_0205_),
    .B2(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0038_));
 sky130_fd_sc_hd__and3_1 _1336_ (.A(net13),
    .B(\UARTReceiver_ins.data[5] ),
    .C(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0211_));
 sky130_fd_sc_hd__o22a_1 _1337_ (.A1(\SRAMController_ins.rx_data_out[5] ),
    .A2(_0204_),
    .B1(_0205_),
    .B2(_0211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0039_));
 sky130_fd_sc_hd__and3_1 _1338_ (.A(net13),
    .B(\UARTReceiver_ins.data[6] ),
    .C(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0212_));
 sky130_fd_sc_hd__o22a_1 _1339_ (.A1(net111),
    .A2(_0204_),
    .B1(_0205_),
    .B2(_0212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0040_));
 sky130_fd_sc_hd__and3_1 _1340_ (.A(net13),
    .B(\UARTReceiver_ins.data[7] ),
    .C(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0213_));
 sky130_fd_sc_hd__o22a_1 _1341_ (.A1(\SRAMController_ins.rx_data_out[7] ),
    .A2(_0204_),
    .B1(_0205_),
    .B2(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0041_));
 sky130_fd_sc_hd__a21boi_1 _1342_ (.A1(\UARTTransmitter_ins.txCounter[0] ),
    .A2(_0423_),
    .B1_N(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0214_));
 sky130_fd_sc_hd__o21a_1 _1343_ (.A1(net109),
    .A2(_0423_),
    .B1(_0214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0042_));
 sky130_fd_sc_hd__and3_1 _1344_ (.A(\UARTTransmitter_ins.txCounter[1] ),
    .B(\UARTTransmitter_ins.txCounter[0] ),
    .C(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0215_));
 sky130_fd_sc_hd__a21o_1 _1345_ (.A1(\UARTTransmitter_ins.txCounter[0] ),
    .A2(_0423_),
    .B1(\UARTTransmitter_ins.txCounter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0216_));
 sky130_fd_sc_hd__and3b_1 _1346_ (.A_N(_0215_),
    .B(_0216_),
    .C(_0429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0217_));
 sky130_fd_sc_hd__clkbuf_1 _1347_ (.A(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _1348_ (.A(\UARTTransmitter_ins.txCounter[2] ),
    .B(_0215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0218_));
 sky130_fd_sc_hd__o21ai_1 _1349_ (.A1(net103),
    .A2(_0215_),
    .B1(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0219_));
 sky130_fd_sc_hd__nor2_1 _1350_ (.A(_0218_),
    .B(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0044_));
 sky130_fd_sc_hd__and3_1 _1351_ (.A(\UARTTransmitter_ins.txCounter[3] ),
    .B(\UARTTransmitter_ins.txCounter[2] ),
    .C(_0215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0220_));
 sky130_fd_sc_hd__o21ai_1 _1352_ (.A1(net95),
    .A2(_0218_),
    .B1(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0221_));
 sky130_fd_sc_hd__nor2_1 _1353_ (.A(_0220_),
    .B(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0045_));
 sky130_fd_sc_hd__and2_1 _1354_ (.A(\UARTTransmitter_ins.txCounter[4] ),
    .B(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0222_));
 sky130_fd_sc_hd__o21ai_1 _1355_ (.A1(net102),
    .A2(_0220_),
    .B1(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0223_));
 sky130_fd_sc_hd__nor2_1 _1356_ (.A(_0222_),
    .B(_0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0046_));
 sky130_fd_sc_hd__and3_1 _1357_ (.A(\UARTTransmitter_ins.txCounter[5] ),
    .B(\UARTTransmitter_ins.txCounter[4] ),
    .C(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0224_));
 sky130_fd_sc_hd__o21ai_1 _1358_ (.A1(net98),
    .A2(_0222_),
    .B1(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0225_));
 sky130_fd_sc_hd__nor2_1 _1359_ (.A(_0224_),
    .B(_0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0047_));
 sky130_fd_sc_hd__and2_1 _1360_ (.A(\UARTTransmitter_ins.txCounter[6] ),
    .B(_0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0226_));
 sky130_fd_sc_hd__o21ai_1 _1361_ (.A1(net114),
    .A2(_0224_),
    .B1(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0227_));
 sky130_fd_sc_hd__nor2_1 _1362_ (.A(_0226_),
    .B(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0048_));
 sky130_fd_sc_hd__o21ai_1 _1363_ (.A1(\UARTTransmitter_ins.txCounter[7] ),
    .A2(_0226_),
    .B1(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0228_));
 sky130_fd_sc_hd__a21oi_1 _1364_ (.A1(net86),
    .A2(_0226_),
    .B1(_0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0049_));
 sky130_fd_sc_hd__and3_1 _1365_ (.A(\UARTTransmitter_ins.txCounter[8] ),
    .B(\UARTTransmitter_ins.txCounter[7] ),
    .C(_0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0229_));
 sky130_fd_sc_hd__a31o_1 _1366_ (.A1(\UARTTransmitter_ins.txCounter[7] ),
    .A2(\UARTTransmitter_ins.txCounter[6] ),
    .A3(_0224_),
    .B1(\UARTTransmitter_ins.txCounter[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0230_));
 sky130_fd_sc_hd__and3b_1 _1367_ (.A_N(_0229_),
    .B(_0429_),
    .C(_0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_1 _1368_ (.A(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _1369_ (.A(\UARTTransmitter_ins.txCounter[9] ),
    .B(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0232_));
 sky130_fd_sc_hd__o21ai_1 _1370_ (.A1(net93),
    .A2(_0229_),
    .B1(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0233_));
 sky130_fd_sc_hd__nor2_1 _1371_ (.A(_0232_),
    .B(_0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0051_));
 sky130_fd_sc_hd__or2_1 _1372_ (.A(\UARTTransmitter_ins.txCounter[10] ),
    .B(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0234_));
 sky130_fd_sc_hd__nand2_1 _1373_ (.A(\UARTTransmitter_ins.txCounter[10] ),
    .B(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0235_));
 sky130_fd_sc_hd__and3_1 _1374_ (.A(_0429_),
    .B(_0234_),
    .C(_0235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0236_));
 sky130_fd_sc_hd__clkbuf_1 _1375_ (.A(_0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0052_));
 sky130_fd_sc_hd__inv_2 _1376_ (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0237_));
 sky130_fd_sc_hd__a21boi_1 _1377_ (.A1(_0237_),
    .A2(_0235_),
    .B1_N(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0053_));
 sky130_fd_sc_hd__a21o_2 _1378_ (.A1(\UARTTransmitter_ins.state[0] ),
    .A2(_0409_),
    .B1(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0238_));
 sky130_fd_sc_hd__a22o_1 _1379_ (.A1(\SRAMController_ins.sram_tmp[0] ),
    .A2(_0413_),
    .B1(_0672_),
    .B2(\SRAMController_ins.sram_tmp[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0239_));
 sky130_fd_sc_hd__a221o_2 _1380_ (.A1(\SRAMController_ins.sram_tmp[16] ),
    .A2(_0673_),
    .B1(_0421_),
    .B2(\SRAMController_ins.sram_tmp[24] ),
    .C1(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0240_));
 sky130_fd_sc_hd__a21oi_4 _1381_ (.A1(\UARTTransmitter_ins.state[0] ),
    .A2(_0409_),
    .B1(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0241_));
 sky130_fd_sc_hd__a21o_1 _1382_ (.A1(net17),
    .A2(_0240_),
    .B1(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0242_));
 sky130_fd_sc_hd__o211a_1 _1383_ (.A1(net73),
    .A2(_0238_),
    .B1(_0242_),
    .C1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0054_));
 sky130_fd_sc_hd__a22o_1 _1384_ (.A1(\SRAMController_ins.sram_tmp[1] ),
    .A2(_0413_),
    .B1(_0672_),
    .B2(\SRAMController_ins.sram_tmp[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0243_));
 sky130_fd_sc_hd__a221o_2 _1385_ (.A1(\SRAMController_ins.sram_tmp[17] ),
    .A2(_0673_),
    .B1(_0421_),
    .B2(\SRAMController_ins.sram_tmp[25] ),
    .C1(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0244_));
 sky130_fd_sc_hd__a21o_1 _1386_ (.A1(\SRAMController_ins.tx_ready ),
    .A2(_0244_),
    .B1(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0245_));
 sky130_fd_sc_hd__o211a_1 _1387_ (.A1(net81),
    .A2(_0238_),
    .B1(_0245_),
    .C1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0055_));
 sky130_fd_sc_hd__a22o_1 _1388_ (.A1(\SRAMController_ins.sram_tmp[2] ),
    .A2(_0413_),
    .B1(_0672_),
    .B2(\SRAMController_ins.sram_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0246_));
 sky130_fd_sc_hd__a221o_2 _1389_ (.A1(\SRAMController_ins.sram_tmp[18] ),
    .A2(_0673_),
    .B1(_0421_),
    .B2(\SRAMController_ins.sram_tmp[26] ),
    .C1(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0247_));
 sky130_fd_sc_hd__a21o_1 _1390_ (.A1(\SRAMController_ins.tx_ready ),
    .A2(_0247_),
    .B1(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0248_));
 sky130_fd_sc_hd__o211a_1 _1391_ (.A1(net79),
    .A2(_0238_),
    .B1(_0248_),
    .C1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0056_));
 sky130_fd_sc_hd__a22o_1 _1392_ (.A1(\SRAMController_ins.sram_tmp[3] ),
    .A2(_0413_),
    .B1(_0672_),
    .B2(\SRAMController_ins.sram_tmp[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0249_));
 sky130_fd_sc_hd__a221o_2 _1393_ (.A1(\SRAMController_ins.sram_tmp[19] ),
    .A2(_0673_),
    .B1(_0421_),
    .B2(\SRAMController_ins.sram_tmp[27] ),
    .C1(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0250_));
 sky130_fd_sc_hd__a21o_1 _1394_ (.A1(\SRAMController_ins.tx_ready ),
    .A2(_0250_),
    .B1(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0251_));
 sky130_fd_sc_hd__o211a_1 _1395_ (.A1(net78),
    .A2(_0238_),
    .B1(_0251_),
    .C1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0057_));
 sky130_fd_sc_hd__a22o_1 _1396_ (.A1(\SRAMController_ins.sram_tmp[4] ),
    .A2(_0413_),
    .B1(_0672_),
    .B2(\SRAMController_ins.sram_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0252_));
 sky130_fd_sc_hd__a221o_2 _1397_ (.A1(\SRAMController_ins.sram_tmp[20] ),
    .A2(_0673_),
    .B1(_0421_),
    .B2(\SRAMController_ins.sram_tmp[28] ),
    .C1(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0253_));
 sky130_fd_sc_hd__a21o_1 _1398_ (.A1(net17),
    .A2(_0253_),
    .B1(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0254_));
 sky130_fd_sc_hd__o211a_1 _1399_ (.A1(net80),
    .A2(_0238_),
    .B1(_0254_),
    .C1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0058_));
 sky130_fd_sc_hd__a22o_1 _1400_ (.A1(\SRAMController_ins.sram_tmp[5] ),
    .A2(_0413_),
    .B1(_0672_),
    .B2(\SRAMController_ins.sram_tmp[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0255_));
 sky130_fd_sc_hd__a221o_2 _1401_ (.A1(\SRAMController_ins.sram_tmp[21] ),
    .A2(_0673_),
    .B1(_0421_),
    .B2(\SRAMController_ins.sram_tmp[29] ),
    .C1(_0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0256_));
 sky130_fd_sc_hd__a21o_1 _1402_ (.A1(net17),
    .A2(_0256_),
    .B1(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0257_));
 sky130_fd_sc_hd__o211a_1 _1403_ (.A1(net74),
    .A2(_0238_),
    .B1(_0257_),
    .C1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0059_));
 sky130_fd_sc_hd__a22o_1 _1404_ (.A1(\SRAMController_ins.sram_tmp[6] ),
    .A2(_0413_),
    .B1(_0672_),
    .B2(\SRAMController_ins.sram_tmp[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0258_));
 sky130_fd_sc_hd__a221o_2 _1405_ (.A1(\SRAMController_ins.sram_tmp[22] ),
    .A2(_0673_),
    .B1(_0421_),
    .B2(\SRAMController_ins.sram_tmp[30] ),
    .C1(_0258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0259_));
 sky130_fd_sc_hd__a21o_1 _1406_ (.A1(net17),
    .A2(_0259_),
    .B1(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0260_));
 sky130_fd_sc_hd__o211a_1 _1407_ (.A1(net82),
    .A2(_0238_),
    .B1(_0260_),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0060_));
 sky130_fd_sc_hd__a22o_1 _1408_ (.A1(\SRAMController_ins.sram_tmp[7] ),
    .A2(_0413_),
    .B1(_0672_),
    .B2(\SRAMController_ins.sram_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0261_));
 sky130_fd_sc_hd__a221o_2 _1409_ (.A1(\SRAMController_ins.sram_tmp[23] ),
    .A2(_0673_),
    .B1(_0421_),
    .B2(\SRAMController_ins.sram_tmp[31] ),
    .C1(_0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0262_));
 sky130_fd_sc_hd__a21o_1 _1410_ (.A1(net17),
    .A2(_0262_),
    .B1(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0263_));
 sky130_fd_sc_hd__o211a_1 _1411_ (.A1(net77),
    .A2(_0238_),
    .B1(_0263_),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0061_));
 sky130_fd_sc_hd__and3_1 _1412_ (.A(\UARTTransmitter_ins.state[1] ),
    .B(_0409_),
    .C(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0264_));
 sky130_fd_sc_hd__o21ai_1 _1413_ (.A1(\UARTTransmitter_ins.state[0] ),
    .A2(\UARTTransmitter_ins.state[1] ),
    .B1(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0265_));
 sky130_fd_sc_hd__mux2_1 _1414_ (.A0(_0264_),
    .A1(_0265_),
    .S(\UARTTransmitter_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0266_));
 sky130_fd_sc_hd__and2_1 _1415_ (.A(net29),
    .B(_0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0267_));
 sky130_fd_sc_hd__clkbuf_1 _1416_ (.A(_0267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0062_));
 sky130_fd_sc_hd__o21ai_1 _1417_ (.A1(\UARTTransmitter_ins.bitIndex[1] ),
    .A2(\UARTTransmitter_ins.bitIndex[0] ),
    .B1(_0264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0268_));
 sky130_fd_sc_hd__o2bb2a_1 _1418_ (.A1_N(\UARTTransmitter_ins.bitIndex[1] ),
    .A2_N(_0265_),
    .B1(_0268_),
    .B2(_0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0269_));
 sky130_fd_sc_hd__nor2_1 _1419_ (.A(_0398_),
    .B(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0063_));
 sky130_fd_sc_hd__or2_1 _1420_ (.A(\UARTTransmitter_ins.bitIndex[2] ),
    .B(_0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0270_));
 sky130_fd_sc_hd__a32o_1 _1421_ (.A1(_0431_),
    .A2(_0264_),
    .A3(_0270_),
    .B1(_0265_),
    .B2(\UARTTransmitter_ins.bitIndex[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0271_));
 sky130_fd_sc_hd__and2_1 _1422_ (.A(net28),
    .B(_0271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0272_));
 sky130_fd_sc_hd__clkbuf_1 _1423_ (.A(_0272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0064_));
 sky130_fd_sc_hd__inv_2 _1424_ (.A(\UARTTransmitter_ins.bitIndex[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0273_));
 sky130_fd_sc_hd__mux4_1 _1425_ (.A0(\UARTTransmitter_ins.data[4] ),
    .A1(\UARTTransmitter_ins.data[5] ),
    .A2(\UARTTransmitter_ins.data[6] ),
    .A3(\UARTTransmitter_ins.data[7] ),
    .S0(\UARTTransmitter_ins.bitIndex[0] ),
    .S1(\UARTTransmitter_ins.bitIndex[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0274_));
 sky130_fd_sc_hd__mux4_1 _1426_ (.A0(\UARTTransmitter_ins.data[0] ),
    .A1(\UARTTransmitter_ins.data[1] ),
    .A2(\UARTTransmitter_ins.data[2] ),
    .A3(\UARTTransmitter_ins.data[3] ),
    .S0(\UARTTransmitter_ins.bitIndex[0] ),
    .S1(\UARTTransmitter_ins.bitIndex[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0275_));
 sky130_fd_sc_hd__or2_1 _1427_ (.A(\UARTTransmitter_ins.bitIndex[2] ),
    .B(_0275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0276_));
 sky130_fd_sc_hd__o211a_1 _1428_ (.A1(_0273_),
    .A2(_0274_),
    .B1(_0276_),
    .C1(\UARTTransmitter_ins.state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0277_));
 sky130_fd_sc_hd__or4b_1 _1429_ (.A(_0398_),
    .B(\UARTTransmitter_ins.state[3] ),
    .C(_0277_),
    .D_N(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0278_));
 sky130_fd_sc_hd__o32a_1 _1430_ (.A1(net75),
    .A2(_0398_),
    .A3(_0428_),
    .B1(_0278_),
    .B2(\UARTTransmitter_ins.state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0065_));
 sky130_fd_sc_hd__a31o_1 _1431_ (.A1(\UARTTransmitter_ins.txCounter[11] ),
    .A2(\UARTTransmitter_ins.state[0] ),
    .A3(_0408_),
    .B1(\SRAMController_ins.tx_ready ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0279_));
 sky130_fd_sc_hd__and3_1 _1432_ (.A(net28),
    .B(_0423_),
    .C(_0279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_1 _1433_ (.A(_0280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1434_ (.A0(\SRAMController_ins.sram_addr_from_dpu[0] ),
    .A1(\SRAMController_ins.rx_data_out[0] ),
    .S(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0281_));
 sky130_fd_sc_hd__clkbuf_1 _1435_ (.A(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1436_ (.A0(\SRAMController_ins.sram_addr_from_dpu[1] ),
    .A1(\SRAMController_ins.rx_data_out[1] ),
    .S(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0282_));
 sky130_fd_sc_hd__clkbuf_1 _1437_ (.A(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1438_ (.A0(\SRAMController_ins.sram_addr_from_dpu[2] ),
    .A1(\SRAMController_ins.rx_data_out[2] ),
    .S(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0283_));
 sky130_fd_sc_hd__clkbuf_1 _1439_ (.A(_0283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(\SRAMController_ins.sram_addr_from_dpu[3] ),
    .A1(\SRAMController_ins.rx_data_out[3] ),
    .S(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0284_));
 sky130_fd_sc_hd__clkbuf_1 _1441_ (.A(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1442_ (.A0(\dpu_ins.cur_cmd[5] ),
    .A1(\SRAMController_ins.rx_data_out[5] ),
    .S(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0285_));
 sky130_fd_sc_hd__clkbuf_1 _1443_ (.A(_0285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(net10),
    .A1(\SRAMController_ins.rx_data_out[6] ),
    .S(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0286_));
 sky130_fd_sc_hd__clkbuf_1 _1445_ (.A(_0286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0072_));
 sky130_fd_sc_hd__and3b_1 _1446_ (.A_N(_0422_),
    .B(_0666_),
    .C(_0200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_8 _1447_ (.A(_0287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0288_));
 sky130_fd_sc_hd__buf_4 _1448_ (.A(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _1449_ (.A0(\SRAMController_ins.sram_tmp[0] ),
    .A1(\SRAMController_ins.sram_data_out[0] ),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0290_));
 sky130_fd_sc_hd__clkbuf_1 _1450_ (.A(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(\SRAMController_ins.sram_tmp[1] ),
    .A1(\SRAMController_ins.sram_data_out[1] ),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _1452_ (.A(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1453_ (.A0(\SRAMController_ins.sram_tmp[2] ),
    .A1(\SRAMController_ins.sram_data_out[2] ),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_1 _1454_ (.A(_0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1455_ (.A0(\SRAMController_ins.sram_tmp[3] ),
    .A1(\SRAMController_ins.sram_data_out[3] ),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _1456_ (.A(_0293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1457_ (.A0(\SRAMController_ins.sram_tmp[4] ),
    .A1(\SRAMController_ins.sram_data_out[4] ),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _1458_ (.A(_0294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1459_ (.A0(\SRAMController_ins.sram_tmp[5] ),
    .A1(\SRAMController_ins.sram_data_out[5] ),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _1460_ (.A(_0295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _1461_ (.A0(\SRAMController_ins.sram_tmp[6] ),
    .A1(\SRAMController_ins.sram_data_out[6] ),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _1462_ (.A(_0296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _1463_ (.A0(\SRAMController_ins.sram_tmp[7] ),
    .A1(\SRAMController_ins.sram_data_out[7] ),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0297_));
 sky130_fd_sc_hd__clkbuf_1 _1464_ (.A(_0297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1465_ (.A0(\SRAMController_ins.sram_tmp[8] ),
    .A1(\SRAMController_ins.sram_data_out[8] ),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_1 _1466_ (.A(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(\SRAMController_ins.sram_tmp[9] ),
    .A1(\SRAMController_ins.sram_data_out[9] ),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _1468_ (.A(_0299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0082_));
 sky130_fd_sc_hd__buf_4 _1469_ (.A(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _1470_ (.A0(\SRAMController_ins.sram_tmp[10] ),
    .A1(\SRAMController_ins.sram_data_out[10] ),
    .S(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _1471_ (.A(_0301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _1472_ (.A0(\SRAMController_ins.sram_tmp[11] ),
    .A1(\SRAMController_ins.sram_data_out[11] ),
    .S(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_1 _1473_ (.A(_0302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _1474_ (.A0(\SRAMController_ins.sram_tmp[12] ),
    .A1(\SRAMController_ins.sram_data_out[12] ),
    .S(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _1475_ (.A(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _1476_ (.A0(\SRAMController_ins.sram_tmp[13] ),
    .A1(\SRAMController_ins.sram_data_out[13] ),
    .S(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_1 _1477_ (.A(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _1478_ (.A0(\SRAMController_ins.sram_tmp[14] ),
    .A1(\SRAMController_ins.sram_data_out[14] ),
    .S(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _1479_ (.A(_0305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _1480_ (.A0(\SRAMController_ins.sram_tmp[15] ),
    .A1(\SRAMController_ins.sram_data_out[15] ),
    .S(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_1 _1481_ (.A(_0306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _1482_ (.A0(\SRAMController_ins.sram_tmp[16] ),
    .A1(\SRAMController_ins.sram_data_out[16] ),
    .S(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_1 _1483_ (.A(_0307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1484_ (.A0(\SRAMController_ins.sram_tmp[17] ),
    .A1(\SRAMController_ins.sram_data_out[17] ),
    .S(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_1 _1485_ (.A(_0308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(\SRAMController_ins.sram_tmp[18] ),
    .A1(\SRAMController_ins.sram_data_out[18] ),
    .S(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_1 _1487_ (.A(_0309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _1488_ (.A0(\SRAMController_ins.sram_tmp[19] ),
    .A1(\SRAMController_ins.sram_data_out[19] ),
    .S(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _1489_ (.A(_0310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_4 _1490_ (.A(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _1491_ (.A0(\SRAMController_ins.sram_tmp[20] ),
    .A1(\SRAMController_ins.sram_data_out[20] ),
    .S(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _1492_ (.A(_0312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1493_ (.A0(\SRAMController_ins.sram_tmp[21] ),
    .A1(\SRAMController_ins.sram_data_out[21] ),
    .S(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _1494_ (.A(_0313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(\SRAMController_ins.sram_tmp[22] ),
    .A1(\SRAMController_ins.sram_data_out[22] ),
    .S(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _1496_ (.A(_0314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _1497_ (.A0(\SRAMController_ins.sram_tmp[23] ),
    .A1(\SRAMController_ins.sram_data_out[23] ),
    .S(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_1 _1498_ (.A(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _1499_ (.A0(\SRAMController_ins.sram_tmp[24] ),
    .A1(\SRAMController_ins.sram_data_out[24] ),
    .S(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_1 _1500_ (.A(_0316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _1501_ (.A0(\SRAMController_ins.sram_tmp[25] ),
    .A1(\SRAMController_ins.sram_data_out[25] ),
    .S(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_1 _1502_ (.A(_0317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _1503_ (.A0(\SRAMController_ins.sram_tmp[26] ),
    .A1(\SRAMController_ins.sram_data_out[26] ),
    .S(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_1 _1504_ (.A(_0318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _1505_ (.A0(\SRAMController_ins.sram_tmp[27] ),
    .A1(\SRAMController_ins.sram_data_out[27] ),
    .S(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _1506_ (.A(_0319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _1507_ (.A0(\SRAMController_ins.sram_tmp[28] ),
    .A1(\SRAMController_ins.sram_data_out[28] ),
    .S(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _1508_ (.A(_0320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1509_ (.A0(\SRAMController_ins.sram_tmp[29] ),
    .A1(\SRAMController_ins.sram_data_out[29] ),
    .S(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _1510_ (.A(_0321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1511_ (.A0(\SRAMController_ins.sram_tmp[30] ),
    .A1(\SRAMController_ins.sram_data_out[30] ),
    .S(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_1 _1512_ (.A(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1513_ (.A0(\SRAMController_ins.sram_tmp[31] ),
    .A1(\SRAMController_ins.sram_data_out[31] ),
    .S(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _1514_ (.A(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0104_));
 sky130_fd_sc_hd__nor2_1 _1515_ (.A(_0687_),
    .B(_0200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0324_));
 sky130_fd_sc_hd__and4b_1 _1516_ (.A_N(\SRAMController_ins.uart_ready ),
    .B(_0677_),
    .C(_0324_),
    .D(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_2 _1517_ (.A(_0325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_4 _1518_ (.A(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _1519_ (.A0(\SRAMController_ins.data_tmp[0] ),
    .A1(\SRAMController_ins.data_tmp[8] ),
    .S(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _1520_ (.A(_0328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1521_ (.A0(\SRAMController_ins.data_tmp[1] ),
    .A1(\SRAMController_ins.data_tmp[9] ),
    .S(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _1522_ (.A(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1523_ (.A0(\SRAMController_ins.data_tmp[2] ),
    .A1(\SRAMController_ins.data_tmp[10] ),
    .S(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _1524_ (.A(_0330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1525_ (.A0(\SRAMController_ins.data_tmp[3] ),
    .A1(\SRAMController_ins.data_tmp[11] ),
    .S(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_1 _1526_ (.A(_0331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1527_ (.A0(\SRAMController_ins.data_tmp[4] ),
    .A1(\SRAMController_ins.data_tmp[12] ),
    .S(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _1528_ (.A(_0332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1529_ (.A0(\SRAMController_ins.data_tmp[5] ),
    .A1(\SRAMController_ins.data_tmp[13] ),
    .S(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_1 _1530_ (.A(_0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _1531_ (.A0(\SRAMController_ins.data_tmp[6] ),
    .A1(\SRAMController_ins.data_tmp[14] ),
    .S(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_1 _1532_ (.A(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _1533_ (.A0(\SRAMController_ins.data_tmp[7] ),
    .A1(\SRAMController_ins.data_tmp[15] ),
    .S(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_1 _1534_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1535_ (.A0(\SRAMController_ins.data_tmp[8] ),
    .A1(\SRAMController_ins.data_tmp[16] ),
    .S(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_1 _1536_ (.A(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1537_ (.A0(\SRAMController_ins.data_tmp[9] ),
    .A1(\SRAMController_ins.data_tmp[17] ),
    .S(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _1538_ (.A(_0337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0114_));
 sky130_fd_sc_hd__buf_4 _1539_ (.A(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _1540_ (.A0(\SRAMController_ins.data_tmp[10] ),
    .A1(\SRAMController_ins.data_tmp[18] ),
    .S(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _1541_ (.A(_0339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _1542_ (.A0(\SRAMController_ins.data_tmp[11] ),
    .A1(\SRAMController_ins.data_tmp[19] ),
    .S(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _1543_ (.A(_0340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _1544_ (.A0(\SRAMController_ins.data_tmp[12] ),
    .A1(\SRAMController_ins.data_tmp[20] ),
    .S(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _1545_ (.A(_0341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1546_ (.A0(\SRAMController_ins.data_tmp[13] ),
    .A1(\SRAMController_ins.data_tmp[21] ),
    .S(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0342_));
 sky130_fd_sc_hd__clkbuf_1 _1547_ (.A(_0342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _1548_ (.A0(\SRAMController_ins.data_tmp[14] ),
    .A1(\SRAMController_ins.data_tmp[22] ),
    .S(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _1549_ (.A(_0343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _1550_ (.A0(\SRAMController_ins.data_tmp[15] ),
    .A1(\SRAMController_ins.data_tmp[23] ),
    .S(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _1551_ (.A(_0344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(\SRAMController_ins.data_tmp[16] ),
    .A1(\SRAMController_ins.data_tmp[24] ),
    .S(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _1553_ (.A(_0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _1554_ (.A0(\SRAMController_ins.data_tmp[17] ),
    .A1(\SRAMController_ins.data_tmp[25] ),
    .S(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_1 _1555_ (.A(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1556_ (.A0(\SRAMController_ins.data_tmp[18] ),
    .A1(\SRAMController_ins.data_tmp[26] ),
    .S(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0347_));
 sky130_fd_sc_hd__clkbuf_1 _1557_ (.A(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1558_ (.A0(\SRAMController_ins.data_tmp[19] ),
    .A1(\SRAMController_ins.data_tmp[27] ),
    .S(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0348_));
 sky130_fd_sc_hd__clkbuf_1 _1559_ (.A(_0348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_8 _1560_ (.A(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _1561_ (.A0(\SRAMController_ins.data_tmp[20] ),
    .A1(\SRAMController_ins.data_tmp[28] ),
    .S(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0350_));
 sky130_fd_sc_hd__clkbuf_1 _1562_ (.A(_0350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _1563_ (.A0(\SRAMController_ins.data_tmp[21] ),
    .A1(\SRAMController_ins.data_tmp[29] ),
    .S(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _1564_ (.A(_0351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1565_ (.A0(\SRAMController_ins.data_tmp[22] ),
    .A1(\SRAMController_ins.data_tmp[30] ),
    .S(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_1 _1566_ (.A(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(\SRAMController_ins.data_tmp[23] ),
    .A1(\SRAMController_ins.data_tmp[31] ),
    .S(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _1568_ (.A(_0353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _1569_ (.A0(\SRAMController_ins.data_tmp[24] ),
    .A1(\SRAMController_ins.rx_data_out[0] ),
    .S(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _1570_ (.A(_0354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _1571_ (.A0(\SRAMController_ins.data_tmp[25] ),
    .A1(\SRAMController_ins.rx_data_out[1] ),
    .S(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _1572_ (.A(_0355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _1573_ (.A0(\SRAMController_ins.data_tmp[26] ),
    .A1(\SRAMController_ins.rx_data_out[2] ),
    .S(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _1574_ (.A(_0356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _1575_ (.A0(\SRAMController_ins.data_tmp[27] ),
    .A1(\SRAMController_ins.rx_data_out[3] ),
    .S(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _1576_ (.A(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _1577_ (.A0(\SRAMController_ins.data_tmp[28] ),
    .A1(\SRAMController_ins.rx_data_out[4] ),
    .S(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0358_));
 sky130_fd_sc_hd__clkbuf_1 _1578_ (.A(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1579_ (.A0(\SRAMController_ins.data_tmp[29] ),
    .A1(\SRAMController_ins.rx_data_out[5] ),
    .S(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _1580_ (.A(_0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _1581_ (.A0(\SRAMController_ins.data_tmp[30] ),
    .A1(\SRAMController_ins.rx_data_out[6] ),
    .S(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _1582_ (.A(_0360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _1583_ (.A0(\SRAMController_ins.data_tmp[31] ),
    .A1(\SRAMController_ins.rx_data_out[7] ),
    .S(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_1 _1584_ (.A(_0361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0136_));
 sky130_fd_sc_hd__nor2_1 _1585_ (.A(net69),
    .B(_0389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0137_));
 sky130_fd_sc_hd__nand2_1 _1586_ (.A(\UARTReceiver_ins.rxCounter[0] ),
    .B(\UARTReceiver_ins.rxCounter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0362_));
 sky130_fd_sc_hd__and3_1 _1587_ (.A(_0382_),
    .B(_0434_),
    .C(_0362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_1 _1588_ (.A(_0363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0138_));
 sky130_fd_sc_hd__and3_1 _1589_ (.A(\UARTReceiver_ins.rxCounter[0] ),
    .B(\UARTReceiver_ins.rxCounter[2] ),
    .C(\UARTReceiver_ins.rxCounter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0364_));
 sky130_fd_sc_hd__a21o_1 _1590_ (.A1(\UARTReceiver_ins.rxCounter[0] ),
    .A2(\UARTReceiver_ins.rxCounter[1] ),
    .B1(\UARTReceiver_ins.rxCounter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0365_));
 sky130_fd_sc_hd__and3b_1 _1591_ (.A_N(_0364_),
    .B(_0365_),
    .C(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _1592_ (.A(_0366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0139_));
 sky130_fd_sc_hd__and2_1 _1593_ (.A(\UARTReceiver_ins.rxCounter[3] ),
    .B(_0364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0367_));
 sky130_fd_sc_hd__or2_1 _1594_ (.A(\UARTReceiver_ins.rxCounter[3] ),
    .B(_0364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0368_));
 sky130_fd_sc_hd__and3b_1 _1595_ (.A_N(_0367_),
    .B(_0368_),
    .C(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _1596_ (.A(_0369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0140_));
 sky130_fd_sc_hd__and3_1 _1597_ (.A(\UARTReceiver_ins.rxCounter[4] ),
    .B(\UARTReceiver_ins.rxCounter[3] ),
    .C(_0364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0370_));
 sky130_fd_sc_hd__o21ai_1 _1598_ (.A1(net105),
    .A2(_0367_),
    .B1(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0371_));
 sky130_fd_sc_hd__nor2_1 _1599_ (.A(_0370_),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0141_));
 sky130_fd_sc_hd__and3_1 _1600_ (.A(\UARTReceiver_ins.rxCounter[5] ),
    .B(\UARTReceiver_ins.rxCounter[4] ),
    .C(_0367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0372_));
 sky130_fd_sc_hd__o21ai_1 _1601_ (.A1(net97),
    .A2(_0370_),
    .B1(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0373_));
 sky130_fd_sc_hd__nor2_1 _1602_ (.A(_0372_),
    .B(_0373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0142_));
 sky130_fd_sc_hd__o21ai_1 _1603_ (.A1(\UARTReceiver_ins.rxCounter[6] ),
    .A2(_0372_),
    .B1(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0374_));
 sky130_fd_sc_hd__a21oi_1 _1604_ (.A1(net106),
    .A2(_0372_),
    .B1(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0143_));
 sky130_fd_sc_hd__a21oi_1 _1605_ (.A1(\UARTReceiver_ins.rxCounter[6] ),
    .A2(_0372_),
    .B1(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0375_));
 sky130_fd_sc_hd__nor2_1 _1606_ (.A(_0389_),
    .B(_0375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0144_));
 sky130_fd_sc_hd__nor2_4 _1607_ (.A(net9),
    .B(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0376_));
 sky130_fd_sc_hd__clkbuf_4 _1608_ (.A(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0377_));
 sky130_fd_sc_hd__a22o_1 _1609_ (.A1(\dpu_ins.data_in[0] ),
    .A2(_0716_),
    .B1(_0377_),
    .B2(\SRAMController_ins.sram_tmp[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0145_));
 sky130_fd_sc_hd__a22o_1 _1610_ (.A1(\dpu_ins.data_in[1] ),
    .A2(_0716_),
    .B1(_0377_),
    .B2(\SRAMController_ins.sram_tmp[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_1 _1611_ (.A1(\dpu_ins.data_in[2] ),
    .A2(_0716_),
    .B1(_0377_),
    .B2(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0147_));
 sky130_fd_sc_hd__a22o_1 _1612_ (.A1(\dpu_ins.data_in[3] ),
    .A2(_0716_),
    .B1(_0377_),
    .B2(\SRAMController_ins.sram_tmp[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0148_));
 sky130_fd_sc_hd__a22o_1 _1613_ (.A1(\dpu_ins.data_in[4] ),
    .A2(_0716_),
    .B1(_0377_),
    .B2(\SRAMController_ins.sram_tmp[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0149_));
 sky130_fd_sc_hd__a22o_1 _1614_ (.A1(\dpu_ins.data_in[5] ),
    .A2(_0716_),
    .B1(_0377_),
    .B2(\SRAMController_ins.sram_tmp[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_1 _1615_ (.A1(\dpu_ins.data_in[6] ),
    .A2(_0716_),
    .B1(_0377_),
    .B2(\SRAMController_ins.sram_tmp[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0151_));
 sky130_fd_sc_hd__a22o_1 _1616_ (.A1(\dpu_ins.data_in[7] ),
    .A2(_0716_),
    .B1(_0377_),
    .B2(\SRAMController_ins.sram_tmp[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0152_));
 sky130_fd_sc_hd__a22o_1 _1617_ (.A1(\dpu_ins.data_in[8] ),
    .A2(_0716_),
    .B1(_0377_),
    .B2(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_4 _1618_ (.A(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0378_));
 sky130_fd_sc_hd__a22o_1 _1619_ (.A1(\dpu_ins.data_in[9] ),
    .A2(_0378_),
    .B1(_0377_),
    .B2(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0154_));
 sky130_fd_sc_hd__buf_2 _1620_ (.A(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0379_));
 sky130_fd_sc_hd__a22o_1 _1621_ (.A1(\dpu_ins.data_in[10] ),
    .A2(_0378_),
    .B1(_0379_),
    .B2(\SRAMController_ins.sram_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0155_));
 sky130_fd_sc_hd__a22o_1 _1622_ (.A1(\dpu_ins.data_in[11] ),
    .A2(_0378_),
    .B1(_0379_),
    .B2(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0156_));
 sky130_fd_sc_hd__a22o_1 _1623_ (.A1(\dpu_ins.data_in[12] ),
    .A2(_0378_),
    .B1(_0379_),
    .B2(\SRAMController_ins.sram_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0157_));
 sky130_fd_sc_hd__a22o_1 _1624_ (.A1(\dpu_ins.data_in[13] ),
    .A2(_0378_),
    .B1(_0379_),
    .B2(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0158_));
 sky130_fd_sc_hd__a22o_1 _1625_ (.A1(\dpu_ins.data_in[14] ),
    .A2(_0378_),
    .B1(_0379_),
    .B2(\SRAMController_ins.sram_tmp[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_1 _1626_ (.A1(\dpu_ins.data_in[15] ),
    .A2(_0378_),
    .B1(_0379_),
    .B2(\SRAMController_ins.sram_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0160_));
 sky130_fd_sc_hd__a22o_1 _1627_ (.A1(\dpu_ins.data_in[16] ),
    .A2(_0378_),
    .B1(_0379_),
    .B2(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0161_));
 sky130_fd_sc_hd__a22o_1 _1628_ (.A1(\dpu_ins.data_in[17] ),
    .A2(_0378_),
    .B1(_0379_),
    .B2(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_1 _1629_ (.A1(\dpu_ins.data_in[18] ),
    .A2(_0378_),
    .B1(_0379_),
    .B2(\SRAMController_ins.sram_tmp[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0163_));
 sky130_fd_sc_hd__clkbuf_4 _1630_ (.A(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0380_));
 sky130_fd_sc_hd__a22o_1 _1631_ (.A1(\dpu_ins.data_in[19] ),
    .A2(_0380_),
    .B1(_0379_),
    .B2(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0164_));
 sky130_fd_sc_hd__buf_2 _1632_ (.A(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0381_));
 sky130_fd_sc_hd__a22o_1 _1633_ (.A1(\dpu_ins.data_in[20] ),
    .A2(_0380_),
    .B1(_0381_),
    .B2(\SRAMController_ins.sram_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0165_));
 sky130_fd_sc_hd__a22o_1 _1634_ (.A1(\dpu_ins.data_in[21] ),
    .A2(_0380_),
    .B1(_0381_),
    .B2(\SRAMController_ins.sram_tmp[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0166_));
 sky130_fd_sc_hd__a22o_1 _1635_ (.A1(\dpu_ins.data_in[22] ),
    .A2(_0380_),
    .B1(_0381_),
    .B2(\SRAMController_ins.sram_tmp[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _1636_ (.A1(\dpu_ins.data_in[23] ),
    .A2(_0380_),
    .B1(_0381_),
    .B2(\SRAMController_ins.sram_tmp[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_1 _1637_ (.A1(\dpu_ins.data_in[24] ),
    .A2(_0380_),
    .B1(_0381_),
    .B2(\SRAMController_ins.sram_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_1 _1638_ (.A1(\dpu_ins.data_in[25] ),
    .A2(_0380_),
    .B1(_0381_),
    .B2(\SRAMController_ins.sram_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0170_));
 sky130_fd_sc_hd__a22o_1 _1639_ (.A1(\dpu_ins.data_in[26] ),
    .A2(_0380_),
    .B1(_0381_),
    .B2(\SRAMController_ins.sram_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0171_));
 sky130_fd_sc_hd__a22o_1 _1640_ (.A1(\dpu_ins.data_in[27] ),
    .A2(_0380_),
    .B1(_0381_),
    .B2(\SRAMController_ins.sram_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0172_));
 sky130_fd_sc_hd__a22o_1 _1641_ (.A1(\dpu_ins.data_in[28] ),
    .A2(_0380_),
    .B1(_0381_),
    .B2(\SRAMController_ins.sram_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0173_));
 sky130_fd_sc_hd__a22o_1 _1642_ (.A1(\dpu_ins.data_in[29] ),
    .A2(_0715_),
    .B1(_0381_),
    .B2(\SRAMController_ins.sram_tmp[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_1 _1643_ (.A1(net118),
    .A2(_0715_),
    .B1(_0376_),
    .B2(\SRAMController_ins.sram_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_1 _1644_ (.A1(\dpu_ins.data_in[31] ),
    .A2(_0715_),
    .B1(_0376_),
    .B2(\SRAMController_ins.sram_tmp[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0176_));
 sky130_fd_sc_hd__dfxtp_1 _1645_ (.CLK(clknet_leaf_2_clk),
    .D(_0008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.out_latched ));
 sky130_fd_sc_hd__dfxtp_1 _1646_ (.CLK(clknet_leaf_0_clk),
    .D(_0009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1647_ (.CLK(clknet_leaf_17_clk),
    .D(_0010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1648_ (.CLK(clknet_leaf_0_clk),
    .D(_0011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1649_ (.CLK(clknet_leaf_17_clk),
    .D(_0012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1650_ (.CLK(clknet_leaf_17_clk),
    .D(_0013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1651_ (.CLK(clknet_leaf_17_clk),
    .D(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1652_ (.CLK(clknet_leaf_0_clk),
    .D(_0015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1653_ (.CLK(clknet_leaf_0_clk),
    .D(_0016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1654_ (.CLK(clknet_leaf_0_clk),
    .D(_0017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.sampleCount[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1655_ (.CLK(clknet_leaf_0_clk),
    .D(_0018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.sampleCount[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1656_ (.CLK(clknet_leaf_1_clk),
    .D(_0019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.sampleCount[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1657_ (.CLK(clknet_leaf_0_clk),
    .D(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.sampleCount[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1658_ (.CLK(clknet_leaf_1_clk),
    .D(_0021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.inputReg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1659_ (.CLK(clknet_leaf_1_clk),
    .D(_0022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.inputReg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1660_ (.CLK(clknet_leaf_1_clk),
    .D(_0023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.inputReg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1661_ (.CLK(clknet_leaf_0_clk),
    .D(_0024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.bitIndex[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1662_ (.CLK(clknet_leaf_0_clk),
    .D(_0025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.bitIndex[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1663_ (.CLK(clknet_leaf_0_clk),
    .D(_0026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.bitIndex[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1664_ (.CLK(clknet_leaf_0_clk),
    .D(_0027_),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.addr_tmp[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1665_ (.CLK(clknet_leaf_0_clk),
    .D(_0028_),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.addr_tmp[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1666_ (.CLK(clknet_leaf_0_clk),
    .D(_0029_),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.addr_tmp[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1667_ (.CLK(clknet_leaf_1_clk),
    .D(_0030_),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.addr_tmp[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1668_ (.CLK(clknet_leaf_2_clk),
    .D(_0031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.overrun ));
 sky130_fd_sc_hd__dfxtp_1 _1669_ (.CLK(clknet_leaf_3_clk),
    .D(_0032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.error ));
 sky130_fd_sc_hd__dfxtp_1 _1670_ (.CLK(clknet_leaf_2_clk),
    .D(_0033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_valid ));
 sky130_fd_sc_hd__dfxtp_1 _1671_ (.CLK(clknet_leaf_18_clk),
    .D(_0034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1672_ (.CLK(clknet_leaf_17_clk),
    .D(_0035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1673_ (.CLK(clknet_leaf_17_clk),
    .D(_0036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1674_ (.CLK(clknet_leaf_17_clk),
    .D(_0037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1675_ (.CLK(clknet_leaf_17_clk),
    .D(_0038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1676_ (.CLK(clknet_leaf_17_clk),
    .D(_0039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1677_ (.CLK(clknet_leaf_18_clk),
    .D(_0040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1678_ (.CLK(clknet_leaf_0_clk),
    .D(_0041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1679_ (.CLK(clknet_leaf_3_clk),
    .D(_0042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1680_ (.CLK(clknet_leaf_3_clk),
    .D(_0043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1681_ (.CLK(clknet_leaf_3_clk),
    .D(_0044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1682_ (.CLK(clknet_leaf_3_clk),
    .D(_0045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1683_ (.CLK(clknet_leaf_3_clk),
    .D(_0046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1684_ (.CLK(clknet_leaf_3_clk),
    .D(_0047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1685_ (.CLK(clknet_leaf_4_clk),
    .D(_0048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1686_ (.CLK(clknet_leaf_4_clk),
    .D(_0049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1687_ (.CLK(clknet_leaf_4_clk),
    .D(_0050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1688_ (.CLK(clknet_leaf_4_clk),
    .D(_0051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1689_ (.CLK(clknet_leaf_4_clk),
    .D(_0052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1690_ (.CLK(clknet_leaf_4_clk),
    .D(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1691_ (.CLK(clknet_leaf_5_clk),
    .D(_0054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1692_ (.CLK(clknet_leaf_5_clk),
    .D(_0055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1693_ (.CLK(clknet_leaf_4_clk),
    .D(_0056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1694_ (.CLK(clknet_leaf_4_clk),
    .D(_0057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1695_ (.CLK(clknet_leaf_4_clk),
    .D(_0058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1696_ (.CLK(clknet_leaf_4_clk),
    .D(_0059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1697_ (.CLK(clknet_leaf_4_clk),
    .D(_0060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1698_ (.CLK(clknet_leaf_4_clk),
    .D(_0061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1699_ (.CLK(clknet_leaf_4_clk),
    .D(_0062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.bitIndex[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1700_ (.CLK(clknet_leaf_4_clk),
    .D(_0063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.bitIndex[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1701_ (.CLK(clknet_leaf_4_clk),
    .D(_0064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.bitIndex[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1702_ (.CLK(clknet_leaf_4_clk),
    .D(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.out ));
 sky130_fd_sc_hd__dfxtp_1 _1703_ (.CLK(clknet_leaf_3_clk),
    .D(_0066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.tx_ready ));
 sky130_fd_sc_hd__dfxtp_2 _1704_ (.CLK(clknet_leaf_3_clk),
    .D(_0004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1705_ (.CLK(clknet_leaf_4_clk),
    .D(_0005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1706_ (.CLK(clknet_leaf_4_clk),
    .D(_0006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1707_ (.CLK(clknet_leaf_4_clk),
    .D(_0007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1708_ (.CLK(clknet_leaf_1_clk),
    .D(_0000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1709_ (.CLK(clknet_leaf_0_clk),
    .D(_0001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1710_ (.CLK(clknet_leaf_1_clk),
    .D(_0002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1711_ (.CLK(clknet_leaf_0_clk),
    .D(_0003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1712_ (.CLK(clknet_leaf_0_clk),
    .D(_0067_),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_addr_from_dpu[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1713_ (.CLK(clknet_leaf_0_clk),
    .D(_0068_),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_addr_from_dpu[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1714_ (.CLK(clknet_leaf_18_clk),
    .D(_0069_),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_addr_from_dpu[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1715_ (.CLK(clknet_leaf_0_clk),
    .D(_0070_),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_addr_from_dpu[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1716_ (.CLK(clknet_leaf_2_clk),
    .D(_0071_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.cur_cmd[5] ));
 sky130_fd_sc_hd__dfrtp_4 _1717_ (.CLK(clknet_leaf_2_clk),
    .D(_0072_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.cur_cmd[6] ));
 sky130_fd_sc_hd__dfrtp_4 _1718_ (.CLK(clknet_leaf_1_clk),
    .D(\SRAMController_ins.nxt_state[0] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.cur_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1719_ (.CLK(clknet_leaf_1_clk),
    .D(\SRAMController_ins.nxt_state[1] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.cur_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1720_ (.CLK(clknet_leaf_2_clk),
    .D(\SRAMController_ins.nxt_state[2] ),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.cur_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1721_ (.CLK(clknet_leaf_2_clk),
    .D(\SRAMController_ins.nxt_state[3] ),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.cur_state[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1722_ (.CLK(clknet_leaf_14_clk),
    .D(_0073_),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1723_ (.CLK(clknet_leaf_13_clk),
    .D(_0074_),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1724_ (.CLK(clknet_leaf_6_clk),
    .D(_0075_),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1725_ (.CLK(clknet_leaf_7_clk),
    .D(_0076_),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1726_ (.CLK(clknet_leaf_13_clk),
    .D(_0077_),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1727_ (.CLK(clknet_leaf_7_clk),
    .D(_0078_),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1728_ (.CLK(clknet_leaf_7_clk),
    .D(_0079_),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1729_ (.CLK(clknet_leaf_7_clk),
    .D(_0080_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1730_ (.CLK(clknet_leaf_6_clk),
    .D(_0081_),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1731_ (.CLK(clknet_leaf_6_clk),
    .D(_0082_),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[9] ));
 sky130_fd_sc_hd__dfrtp_4 _1732_ (.CLK(clknet_leaf_13_clk),
    .D(_0083_),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1733_ (.CLK(clknet_leaf_7_clk),
    .D(_0084_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[11] ));
 sky130_fd_sc_hd__dfrtp_4 _1734_ (.CLK(clknet_leaf_13_clk),
    .D(_0085_),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1735_ (.CLK(clknet_leaf_7_clk),
    .D(_0086_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[13] ));
 sky130_fd_sc_hd__dfrtp_4 _1736_ (.CLK(clknet_leaf_13_clk),
    .D(_0087_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[14] ));
 sky130_fd_sc_hd__dfrtp_4 _1737_ (.CLK(clknet_leaf_13_clk),
    .D(_0088_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1738_ (.CLK(clknet_leaf_7_clk),
    .D(_0089_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1739_ (.CLK(clknet_leaf_8_clk),
    .D(_0090_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[17] ));
 sky130_fd_sc_hd__dfrtp_4 _1740_ (.CLK(clknet_leaf_13_clk),
    .D(_0091_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1741_ (.CLK(clknet_leaf_8_clk),
    .D(_0092_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[19] ));
 sky130_fd_sc_hd__dfrtp_4 _1742_ (.CLK(clknet_leaf_11_clk),
    .D(_0093_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[20] ));
 sky130_fd_sc_hd__dfrtp_4 _1743_ (.CLK(clknet_leaf_11_clk),
    .D(_0094_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[21] ));
 sky130_fd_sc_hd__dfrtp_4 _1744_ (.CLK(clknet_leaf_12_clk),
    .D(_0095_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[22] ));
 sky130_fd_sc_hd__dfrtp_4 _1745_ (.CLK(clknet_leaf_12_clk),
    .D(_0096_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[23] ));
 sky130_fd_sc_hd__dfrtp_4 _1746_ (.CLK(clknet_leaf_11_clk),
    .D(_0097_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[24] ));
 sky130_fd_sc_hd__dfrtp_4 _1747_ (.CLK(clknet_leaf_11_clk),
    .D(_0098_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[25] ));
 sky130_fd_sc_hd__dfrtp_4 _1748_ (.CLK(clknet_leaf_11_clk),
    .D(_0099_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[26] ));
 sky130_fd_sc_hd__dfrtp_4 _1749_ (.CLK(clknet_leaf_11_clk),
    .D(_0100_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[27] ));
 sky130_fd_sc_hd__dfrtp_4 _1750_ (.CLK(clknet_leaf_11_clk),
    .D(_0101_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[28] ));
 sky130_fd_sc_hd__dfrtp_4 _1751_ (.CLK(clknet_leaf_11_clk),
    .D(_0102_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1752_ (.CLK(clknet_leaf_8_clk),
    .D(_0103_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1753_ (.CLK(clknet_leaf_8_clk),
    .D(_0104_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1754_ (.CLK(clknet_leaf_15_clk),
    .D(_0105_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1755_ (.CLK(clknet_leaf_15_clk),
    .D(_0106_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1756_ (.CLK(clknet_leaf_15_clk),
    .D(_0107_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1757_ (.CLK(clknet_leaf_15_clk),
    .D(_0108_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1758_ (.CLK(clknet_leaf_15_clk),
    .D(_0109_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1759_ (.CLK(clknet_leaf_14_clk),
    .D(_0110_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1760_ (.CLK(clknet_leaf_14_clk),
    .D(_0111_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1761_ (.CLK(clknet_leaf_14_clk),
    .D(_0112_),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1762_ (.CLK(clknet_leaf_15_clk),
    .D(_0113_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1763_ (.CLK(clknet_leaf_15_clk),
    .D(_0114_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[9] ));
 sky130_fd_sc_hd__dfrtp_2 _1764_ (.CLK(clknet_leaf_15_clk),
    .D(_0115_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1765_ (.CLK(clknet_leaf_14_clk),
    .D(_0116_),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1766_ (.CLK(clknet_leaf_13_clk),
    .D(_0117_),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[12] ));
 sky130_fd_sc_hd__dfrtp_4 _1767_ (.CLK(clknet_leaf_12_clk),
    .D(_0118_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[13] ));
 sky130_fd_sc_hd__dfrtp_4 _1768_ (.CLK(clknet_leaf_12_clk),
    .D(_0119_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[14] ));
 sky130_fd_sc_hd__dfrtp_2 _1769_ (.CLK(clknet_leaf_12_clk),
    .D(_0120_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[15] ));
 sky130_fd_sc_hd__dfrtp_4 _1770_ (.CLK(clknet_leaf_15_clk),
    .D(_0121_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[16] ));
 sky130_fd_sc_hd__dfrtp_4 _1771_ (.CLK(clknet_leaf_15_clk),
    .D(_0122_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[17] ));
 sky130_fd_sc_hd__dfrtp_2 _1772_ (.CLK(clknet_leaf_15_clk),
    .D(_0123_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1773_ (.CLK(clknet_leaf_14_clk),
    .D(_0124_),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[19] ));
 sky130_fd_sc_hd__dfrtp_4 _1774_ (.CLK(clknet_leaf_12_clk),
    .D(_0125_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1775_ (.CLK(clknet_leaf_12_clk),
    .D(_0126_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1776_ (.CLK(clknet_leaf_12_clk),
    .D(_0127_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1777_ (.CLK(clknet_leaf_12_clk),
    .D(_0128_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[23] ));
 sky130_fd_sc_hd__dfrtp_4 _1778_ (.CLK(clknet_leaf_16_clk),
    .D(_0129_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[24] ));
 sky130_fd_sc_hd__dfrtp_4 _1779_ (.CLK(clknet_leaf_16_clk),
    .D(_0130_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[25] ));
 sky130_fd_sc_hd__dfrtp_4 _1780_ (.CLK(clknet_leaf_16_clk),
    .D(_0131_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[26] ));
 sky130_fd_sc_hd__dfrtp_4 _1781_ (.CLK(clknet_leaf_16_clk),
    .D(_0132_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[27] ));
 sky130_fd_sc_hd__dfrtp_4 _1782_ (.CLK(clknet_leaf_15_clk),
    .D(_0133_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[28] ));
 sky130_fd_sc_hd__dfrtp_4 _1783_ (.CLK(clknet_leaf_16_clk),
    .D(_0134_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[29] ));
 sky130_fd_sc_hd__dfrtp_4 _1784_ (.CLK(clknet_leaf_17_clk),
    .D(_0135_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[30] ));
 sky130_fd_sc_hd__dfrtp_4 _1785_ (.CLK(clknet_leaf_17_clk),
    .D(_0136_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[31] ));
 sky130_fd_sc_hd__dfxtp_1 _1786_ (.CLK(clknet_leaf_1_clk),
    .D(_0137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1787_ (.CLK(clknet_leaf_1_clk),
    .D(_0138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1788_ (.CLK(clknet_leaf_3_clk),
    .D(_0139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1789_ (.CLK(clknet_leaf_3_clk),
    .D(_0140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1790_ (.CLK(clknet_leaf_3_clk),
    .D(_0141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1791_ (.CLK(clknet_leaf_3_clk),
    .D(_0142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1792_ (.CLK(clknet_leaf_3_clk),
    .D(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1793_ (.CLK(clknet_leaf_2_clk),
    .D(_0144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1794_ (.CLK(clknet_leaf_17_clk),
    .D(\dpu_ins.data_out[0] ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1795_ (.CLK(clknet_leaf_5_clk),
    .D(\dpu_ins.data_out[1] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1796_ (.CLK(clknet_leaf_5_clk),
    .D(\dpu_ins.data_out[2] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1797_ (.CLK(clknet_leaf_6_clk),
    .D(\dpu_ins.data_out[3] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1798_ (.CLK(clknet_leaf_5_clk),
    .D(\dpu_ins.data_out[4] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1799_ (.CLK(clknet_leaf_6_clk),
    .D(\dpu_ins.data_out[5] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[5] ));
 sky130_fd_sc_hd__dfrtp_2 _1800_ (.CLK(clknet_leaf_6_clk),
    .D(\dpu_ins.data_out[6] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[6] ));
 sky130_fd_sc_hd__dfrtp_2 _1801_ (.CLK(clknet_leaf_6_clk),
    .D(\dpu_ins.data_out[7] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[7] ));
 sky130_fd_sc_hd__dfrtp_2 _1802_ (.CLK(clknet_leaf_6_clk),
    .D(\dpu_ins.data_out[8] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[8] ));
 sky130_fd_sc_hd__dfrtp_2 _1803_ (.CLK(clknet_leaf_6_clk),
    .D(\dpu_ins.data_out[9] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[9] ));
 sky130_fd_sc_hd__dfrtp_2 _1804_ (.CLK(clknet_leaf_6_clk),
    .D(\dpu_ins.data_out[10] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[10] ));
 sky130_fd_sc_hd__dfrtp_2 _1805_ (.CLK(clknet_leaf_6_clk),
    .D(\dpu_ins.data_out[11] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[11] ));
 sky130_fd_sc_hd__dfrtp_2 _1806_ (.CLK(clknet_leaf_6_clk),
    .D(\dpu_ins.data_out[12] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[12] ));
 sky130_fd_sc_hd__dfrtp_2 _1807_ (.CLK(clknet_leaf_7_clk),
    .D(\dpu_ins.data_out[13] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[13] ));
 sky130_fd_sc_hd__dfrtp_2 _1808_ (.CLK(clknet_leaf_7_clk),
    .D(\dpu_ins.data_out[14] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[14] ));
 sky130_fd_sc_hd__dfrtp_2 _1809_ (.CLK(clknet_leaf_7_clk),
    .D(\dpu_ins.data_out[15] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[15] ));
 sky130_fd_sc_hd__dfrtp_4 _1810_ (.CLK(clknet_leaf_8_clk),
    .D(\dpu_ins.data_out[16] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[16] ));
 sky130_fd_sc_hd__dfrtp_2 _1811_ (.CLK(clknet_leaf_8_clk),
    .D(\dpu_ins.data_out[17] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[17] ));
 sky130_fd_sc_hd__dfrtp_4 _1812_ (.CLK(clknet_leaf_8_clk),
    .D(\dpu_ins.data_out[18] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[18] ));
 sky130_fd_sc_hd__dfrtp_4 _1813_ (.CLK(clknet_leaf_8_clk),
    .D(\dpu_ins.data_out[19] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[19] ));
 sky130_fd_sc_hd__dfrtp_2 _1814_ (.CLK(clknet_leaf_8_clk),
    .D(\dpu_ins.data_out[20] ),
    .RESET_B(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[20] ));
 sky130_fd_sc_hd__dfrtp_2 _1815_ (.CLK(clknet_leaf_8_clk),
    .D(\dpu_ins.data_out[21] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[21] ));
 sky130_fd_sc_hd__dfrtp_2 _1816_ (.CLK(clknet_leaf_9_clk),
    .D(\dpu_ins.data_out[22] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[22] ));
 sky130_fd_sc_hd__dfrtp_2 _1817_ (.CLK(clknet_leaf_9_clk),
    .D(\dpu_ins.data_out[23] ),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[23] ));
 sky130_fd_sc_hd__dfrtp_4 _1818_ (.CLK(clknet_leaf_9_clk),
    .D(\dpu_ins.data_out[24] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[24] ));
 sky130_fd_sc_hd__dfrtp_4 _1819_ (.CLK(clknet_leaf_9_clk),
    .D(\dpu_ins.data_out[25] ),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[25] ));
 sky130_fd_sc_hd__dfrtp_4 _1820_ (.CLK(clknet_leaf_9_clk),
    .D(\dpu_ins.data_out[26] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[26] ));
 sky130_fd_sc_hd__dfrtp_4 _1821_ (.CLK(clknet_leaf_9_clk),
    .D(\dpu_ins.data_out[27] ),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[27] ));
 sky130_fd_sc_hd__dfrtp_4 _1822_ (.CLK(clknet_leaf_9_clk),
    .D(\dpu_ins.data_out[28] ),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[28] ));
 sky130_fd_sc_hd__dfrtp_4 _1823_ (.CLK(clknet_leaf_10_clk),
    .D(\dpu_ins.data_out[29] ),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[29] ));
 sky130_fd_sc_hd__dfrtp_4 _1824_ (.CLK(clknet_leaf_9_clk),
    .D(\dpu_ins.data_out[30] ),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[30] ));
 sky130_fd_sc_hd__dfrtp_4 _1825_ (.CLK(clknet_leaf_9_clk),
    .D(\dpu_ins.data_out[31] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_data_from_dpu[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1826_ (.CLK(clknet_leaf_2_clk),
    .D(\dpu_ins.nxt_state[0] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.cur_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1827_ (.CLK(clknet_leaf_2_clk),
    .D(\dpu_ins.nxt_state[1] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.cur_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1828_ (.CLK(clknet_leaf_5_clk),
    .D(_0145_),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1829_ (.CLK(clknet_leaf_5_clk),
    .D(_0146_),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1830_ (.CLK(clknet_leaf_6_clk),
    .D(_0147_),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1831_ (.CLK(clknet_leaf_5_clk),
    .D(_0148_),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1832_ (.CLK(clknet_leaf_6_clk),
    .D(_0149_),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1833_ (.CLK(clknet_leaf_5_clk),
    .D(_0150_),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[5] ));
 sky130_fd_sc_hd__dfrtp_2 _1834_ (.CLK(clknet_leaf_6_clk),
    .D(_0151_),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[6] ));
 sky130_fd_sc_hd__dfrtp_2 _1835_ (.CLK(clknet_leaf_6_clk),
    .D(_0152_),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[7] ));
 sky130_fd_sc_hd__dfrtp_2 _1836_ (.CLK(clknet_leaf_6_clk),
    .D(_0153_),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[8] ));
 sky130_fd_sc_hd__dfrtp_2 _1837_ (.CLK(clknet_leaf_6_clk),
    .D(_0154_),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[9] ));
 sky130_fd_sc_hd__dfrtp_2 _1838_ (.CLK(clknet_leaf_7_clk),
    .D(_0155_),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[10] ));
 sky130_fd_sc_hd__dfrtp_2 _1839_ (.CLK(clknet_leaf_7_clk),
    .D(_0156_),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[11] ));
 sky130_fd_sc_hd__dfrtp_2 _1840_ (.CLK(clknet_leaf_7_clk),
    .D(_0157_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[12] ));
 sky130_fd_sc_hd__dfrtp_2 _1841_ (.CLK(clknet_leaf_7_clk),
    .D(_0158_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[13] ));
 sky130_fd_sc_hd__dfrtp_2 _1842_ (.CLK(clknet_leaf_7_clk),
    .D(_0159_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[14] ));
 sky130_fd_sc_hd__dfrtp_2 _1843_ (.CLK(clknet_leaf_7_clk),
    .D(_0160_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[15] ));
 sky130_fd_sc_hd__dfrtp_2 _1844_ (.CLK(clknet_leaf_8_clk),
    .D(_0161_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[16] ));
 sky130_fd_sc_hd__dfrtp_2 _1845_ (.CLK(clknet_leaf_8_clk),
    .D(_0162_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1846_ (.CLK(clknet_leaf_8_clk),
    .D(_0163_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1847_ (.CLK(clknet_leaf_8_clk),
    .D(_0164_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[19] ));
 sky130_fd_sc_hd__dfrtp_4 _1848_ (.CLK(clknet_leaf_10_clk),
    .D(_0165_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[20] ));
 sky130_fd_sc_hd__dfrtp_4 _1849_ (.CLK(clknet_leaf_10_clk),
    .D(_0166_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1850_ (.CLK(clknet_leaf_9_clk),
    .D(_0167_),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[22] ));
 sky130_fd_sc_hd__dfrtp_2 _1851_ (.CLK(clknet_leaf_9_clk),
    .D(_0168_),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[23] ));
 sky130_fd_sc_hd__dfrtp_2 _1852_ (.CLK(clknet_leaf_9_clk),
    .D(_0169_),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[24] ));
 sky130_fd_sc_hd__dfrtp_1 _1853_ (.CLK(clknet_leaf_9_clk),
    .D(_0170_),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[25] ));
 sky130_fd_sc_hd__dfrtp_2 _1854_ (.CLK(clknet_leaf_10_clk),
    .D(_0171_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[26] ));
 sky130_fd_sc_hd__dfrtp_2 _1855_ (.CLK(clknet_leaf_10_clk),
    .D(_0172_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[27] ));
 sky130_fd_sc_hd__dfrtp_1 _1856_ (.CLK(clknet_leaf_10_clk),
    .D(_0173_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1857_ (.CLK(clknet_leaf_9_clk),
    .D(_0174_),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[29] ));
 sky130_fd_sc_hd__dfrtp_2 _1858_ (.CLK(clknet_leaf_9_clk),
    .D(_0175_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1859_ (.CLK(clknet_leaf_9_clk),
    .D(_0176_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\dpu_ins.data_in[31] ));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .HI(net67));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__conb_1 sram_ins_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net43));
 sky130_fd_sc_hd__conb_1 sram_ins_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net44));
 sky130_fd_sc_hd__conb_1 sram_ins_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net45));
 sky130_fd_sc_hd__conb_1 sram_ins_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net46));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net47));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net48));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net49));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net50));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net51));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net52));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net53));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net54));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net55));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net56));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net57));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net58));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net59));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net60));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net61));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net62));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net63));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net64));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net65));
 sky130_fd_sc_hd__conb_1 sram_ins_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .HI(net66));
 sky130_fd_sc_hd__buf_2 _1886_ (.A(\UARTTransmitter_ins.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__clkbuf_4 _1887_ (.A(\SRAMController_ins.uart_ready ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__clkbuf_4 _1888_ (.A(\UARTReceiver_ins.overrun ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__clkbuf_4 _1889_ (.A(\UARTReceiver_ins.error ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(uo_out[7]));
 myconfig_sky_dual sram_ins (.csb0(\SRAMController_ins.csb_n ),
    .csb1(net66),
    .web0(\SRAMController_ins.we_n ),
    .clk0(clknet_leaf_15_clk),
    .clk1(net46),
    .vccd1(VDPWR),
    .vssd1(VGND),
    .addr0({\SRAMController_ins.addr[3] ,
    \SRAMController_ins.addr[2] ,
    \SRAMController_ins.addr[1] ,
    \SRAMController_ins.addr[0] }),
    .addr1({net45,
    net44,
    net43,
    net42}),
    .din0({\SRAMController_ins.sram_data_in[31] ,
    \SRAMController_ins.sram_data_in[30] ,
    \SRAMController_ins.sram_data_in[29] ,
    \SRAMController_ins.sram_data_in[28] ,
    \SRAMController_ins.sram_data_in[27] ,
    \SRAMController_ins.sram_data_in[26] ,
    \SRAMController_ins.sram_data_in[25] ,
    \SRAMController_ins.sram_data_in[24] ,
    \SRAMController_ins.sram_data_in[23] ,
    \SRAMController_ins.sram_data_in[22] ,
    \SRAMController_ins.sram_data_in[21] ,
    \SRAMController_ins.sram_data_in[20] ,
    \SRAMController_ins.sram_data_in[19] ,
    \SRAMController_ins.sram_data_in[18] ,
    \SRAMController_ins.sram_data_in[17] ,
    \SRAMController_ins.sram_data_in[16] ,
    \SRAMController_ins.sram_data_in[15] ,
    \SRAMController_ins.sram_data_in[14] ,
    \SRAMController_ins.sram_data_in[13] ,
    \SRAMController_ins.sram_data_in[12] ,
    \SRAMController_ins.sram_data_in[11] ,
    \SRAMController_ins.sram_data_in[10] ,
    \SRAMController_ins.sram_data_in[9] ,
    \SRAMController_ins.sram_data_in[8] ,
    \SRAMController_ins.sram_data_in[7] ,
    \SRAMController_ins.sram_data_in[6] ,
    \SRAMController_ins.sram_data_in[5] ,
    \SRAMController_ins.sram_data_in[4] ,
    \SRAMController_ins.sram_data_in[3] ,
    \SRAMController_ins.sram_data_in[2] ,
    \SRAMController_ins.sram_data_in[1] ,
    \SRAMController_ins.sram_data_in[0] }),
    .dout0({\SRAMController_ins.sram_data_out[31] ,
    \SRAMController_ins.sram_data_out[30] ,
    \SRAMController_ins.sram_data_out[29] ,
    \SRAMController_ins.sram_data_out[28] ,
    \SRAMController_ins.sram_data_out[27] ,
    \SRAMController_ins.sram_data_out[26] ,
    \SRAMController_ins.sram_data_out[25] ,
    \SRAMController_ins.sram_data_out[24] ,
    \SRAMController_ins.sram_data_out[23] ,
    \SRAMController_ins.sram_data_out[22] ,
    \SRAMController_ins.sram_data_out[21] ,
    \SRAMController_ins.sram_data_out[20] ,
    \SRAMController_ins.sram_data_out[19] ,
    \SRAMController_ins.sram_data_out[18] ,
    \SRAMController_ins.sram_data_out[17] ,
    \SRAMController_ins.sram_data_out[16] ,
    \SRAMController_ins.sram_data_out[15] ,
    \SRAMController_ins.sram_data_out[14] ,
    \SRAMController_ins.sram_data_out[13] ,
    \SRAMController_ins.sram_data_out[12] ,
    \SRAMController_ins.sram_data_out[11] ,
    \SRAMController_ins.sram_data_out[10] ,
    \SRAMController_ins.sram_data_out[9] ,
    \SRAMController_ins.sram_data_out[8] ,
    \SRAMController_ins.sram_data_out[7] ,
    \SRAMController_ins.sram_data_out[6] ,
    \SRAMController_ins.sram_data_out[5] ,
    \SRAMController_ins.sram_data_out[4] ,
    \SRAMController_ins.sram_data_out[3] ,
    \SRAMController_ins.sram_data_out[2] ,
    \SRAMController_ins.sram_data_out[1] ,
    \SRAMController_ins.sram_data_out[0] }),
    .dout1({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_2_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_2_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_2_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_2_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_2_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_2_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_2_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_1_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_1_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_1_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_1_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_1_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_1_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_1_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_2_Left_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_2_Left_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_2_Left_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_2_Left_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_2_Left_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_2_Left_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_2_Left_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Left_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Left_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_1_Right_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_1_Right_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_1_Right_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_1_Right_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_1_Right_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_1_Right_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Right_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Right_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Right_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Right_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Right_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Right_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Right_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Right_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Right_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Right_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Right_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Right_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Right_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Right_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Right_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Right_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Right_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Right_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Right_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Right_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Right_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Right_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Right_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Right_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Right_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Right_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Right_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Right_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Right_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Right_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Right_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Right_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Right_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Right_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Right_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Right_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Right_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Right_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Right_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Right_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Right_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Right_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Right_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Right_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Right_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Right_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Right_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Right_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Right_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Right_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Right_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Right_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Right_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Right_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Right_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Right_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Right_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Right_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Right_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Right_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Right_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Right_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_1_Right_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_300 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_301 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_302 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_303 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_304 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_305 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_306 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_307 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_308 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_309 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_310 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_311 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_312 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_313 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_314 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_315 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_316 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_317 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_318 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_319 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_320 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_321 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_322 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_323 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_324 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_325 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_326 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_327 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_328 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_329 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_330 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_331 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_332 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_333 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_334 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_335 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_336 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_337 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_338 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_339 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_340 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_341 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_342 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_343 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_344 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_345 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_346 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_347 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_348 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_349 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_350 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_351 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_352 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_353 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_354 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_355 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_356 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_357 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_358 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_359 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_360 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_361 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_362 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_363 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_364 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_365 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_366 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_367 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_368 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_369 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_370 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_371 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_372 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_373 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_374 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_375 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_376 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_377 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_378 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_379 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_380 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_381 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_382 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_383 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_384 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_385 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_386 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_387 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_388 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_389 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_390 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_391 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_392 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_393 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_394 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1_395 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1_396 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1_397 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1_398 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1_399 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1_400 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1_401 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1_402 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1_403 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1_404 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1_405 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1_406 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1_407 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1_408 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1_409 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1_410 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1_411 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1_412 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_413 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_414 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_415 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_416 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_417 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_418 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_419 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_420 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_421 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_422 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_423 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_424 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_425 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_426 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_427 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_428 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_429 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_430 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_431 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_432 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_433 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_434 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_435 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_436 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_437 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_438 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_439 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_440 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_441 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_442 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_443 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_444 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_445 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_446 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_447 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_448 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_449 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_450 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_451 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_452 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_453 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_454 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_455 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_456 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_457 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_458 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_459 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_460 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_461 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_462 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_463 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_464 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_465 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_466 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_467 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_468 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_469 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_470 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_471 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_472 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_473 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_474 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_475 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_476 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_477 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_478 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_479 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_480 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_481 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_482 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_483 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_484 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_485 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_486 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_487 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_488 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_489 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_490 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_491 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_492 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_493 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_494 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_495 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_496 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_497 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_498 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_499 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_500 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_501 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_502 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_503 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_504 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_505 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_506 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_507 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_508 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_509 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_510 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_511 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_512 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_513 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_514 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_515 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_516 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_517 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_518 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_519 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_520 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_521 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_522 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_523 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_524 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_525 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_526 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_527 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_528 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_529 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_530 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_531 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_532 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_533 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_534 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_535 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_536 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_537 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_538 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_539 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_540 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_541 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_542 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_543 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_544 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_545 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_546 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_547 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_548 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_549 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_550 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_551 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_552 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_553 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_554 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_555 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_556 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_557 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_558 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_559 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_560 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_561 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_562 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_563 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_564 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_565 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_566 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_567 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_568 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_569 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_570 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_571 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_572 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_573 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_574 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_575 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_576 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_577 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_578 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_579 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_580 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_581 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_582 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_583 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_584 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_585 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_586 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_587 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_588 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_589 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_590 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_591 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_592 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1_593 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1_594 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1_595 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1_596 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1_597 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1_598 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_599 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_600 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_601 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_602 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_603 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_604 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_605 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_606 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_607 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_608 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_609 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_610 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_611 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_612 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_613 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_614 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_615 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_616 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_617 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_618 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_619 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_620 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_621 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_622 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_623 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_624 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_625 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_626 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_627 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_628 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_629 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_630 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_631 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_632 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_633 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_634 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_635 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_636 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_637 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_638 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_639 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_640 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_641 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_642 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_643 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_644 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_645 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_646 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_647 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_648 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_649 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_650 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_651 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_652 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_653 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_654 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_655 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_656 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_657 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_658 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_659 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_660 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_661 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_662 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_663 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_664 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_665 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_666 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_667 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_668 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_669 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_670 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_671 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_672 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_673 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_674 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_675 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_676 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_677 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_678 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_679 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_680 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_681 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_682 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_683 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_684 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_685 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_686 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_687 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_688 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_689 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_690 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_691 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_692 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_693 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_694 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_695 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_696 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_697 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_698 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_699 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_700 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_701 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_702 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_703 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_704 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_705 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_706 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_707 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_708 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_709 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_710 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_711 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_712 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_713 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_714 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_715 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_716 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_717 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_718 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_719 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_720 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_721 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_722 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_723 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_724 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_725 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_726 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_727 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_728 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_729 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_730 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_731 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_732 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_733 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_734 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_735 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_736 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_737 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_738 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_739 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_740 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_741 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_742 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_743 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_744 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_745 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_746 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_747 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_748 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_749 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_750 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_751 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_752 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_753 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_754 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_755 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_756 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_757 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_758 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_759 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_760 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_761 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_762 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_763 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_764 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_765 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_766 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_767 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_768 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_769 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_770 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_771 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_772 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_773 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_774 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_775 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_776 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_777 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_778 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_779 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_780 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_781 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_782 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_783 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_784 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_785 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_786 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_787 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_788 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_789 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_790 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_791 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_792 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_793 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_794 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_795 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_796 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_797 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_798 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_799 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_800 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_801 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_802 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_803 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_804 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_805 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_806 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_807 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1_808 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1_809 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1_810 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_2_811 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_2_812 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_2_813 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_2_814 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_2_815 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_2_816 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_2_817 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_818 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_819 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_820 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_821 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_822 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_823 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_824 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_825 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_826 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_827 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_828 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_829 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_830 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_831 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_832 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_833 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_834 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_835 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_836 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_837 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_838 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_839 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_840 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_841 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_842 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_843 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_844 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_845 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_846 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_847 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_848 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_849 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_850 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_851 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_852 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_853 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_854 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_855 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_856 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_857 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_858 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_859 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_860 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_861 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_862 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_863 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_864 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_865 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_866 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_867 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_868 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_869 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_870 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_871 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_872 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_873 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_874 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_875 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_876 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_877 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_878 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2_879 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__buf_2 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 wire3 (.A(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 max_cap4 (.A(_0612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 max_cap5 (.A(_0693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net5));
 sky130_fd_sc_hd__buf_1 max_cap6 (.A(_0438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 fanout7 (.A(\SRAMController_ins.cur_state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 fanout9 (.A(\SRAMController_ins.cur_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 fanout11 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_4 fanout12 (.A(\dpu_ins.cur_cmd[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(\UARTReceiver_ins.state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 fanout14 (.A(\UARTReceiver_ins.state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net14));
 sky130_fd_sc_hd__buf_2 fanout15 (.A(\UARTReceiver_ins.state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net15));
 sky130_fd_sc_hd__buf_2 fanout16 (.A(\UARTReceiver_ins.state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(\SRAMController_ins.tx_ready ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(\SRAMController_ins.rx_valid ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 fanout19 (.A(\UARTReceiver_ins.bitIndex[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 fanout20 (.A(\UARTReceiver_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 fanout26 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net32));
 sky130_fd_sc_hd__buf_4 fanout33 (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_8 fanout37 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net40));
 sky130_fd_sc_hd__buf_4 fanout41 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net41));
 sky130_fd_sc_hd__conb_1 sram_ins_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net42));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload0 (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload1 (.A(clknet_leaf_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_leaf_1_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_8 clkload3 (.A(clknet_leaf_2_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload4 (.A(clknet_leaf_3_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_8 clkload5 (.A(clknet_leaf_5_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload6 (.A(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_12 clkload7 (.A(clknet_leaf_14_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_leaf_15_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_12 clkload9 (.A(clknet_leaf_16_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_6 clkload10 (.A(clknet_leaf_17_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_12 clkload11 (.A(clknet_leaf_18_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkbuf_8 clkload12 (.A(clknet_leaf_8_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload13 (.A(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_8 clkload14 (.A(clknet_leaf_10_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_6 clkload15 (.A(clknet_leaf_11_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_6 clkload16 (.A(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_6 clkload17 (.A(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\UARTTransmitter_ins.state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\UARTReceiver_ins.rxCounter[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\UARTTransmitter_ins.txCounter[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\UARTTransmitter_ins.state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\UARTTransmitter_ins.data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\UARTTransmitter_ins.data[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\UARTTransmitter_ins.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\UARTTransmitter_ins.data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\UARTTransmitter_ins.data[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\UARTTransmitter_ins.data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\UARTTransmitter_ins.data[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\UARTTransmitter_ins.data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\UARTTransmitter_ins.data[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\UARTReceiver_ins.data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\UARTReceiver_ins.sampleCount[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\UARTTransmitter_ins.txCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\UARTReceiver_ins.inputReg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\UARTTransmitter_ins.state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\SRAMController_ins.sram_tmp[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\UARTReceiver_ins.inputReg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\SRAMController_ins.sram_tmp[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\SRAMController_ins.sram_tmp[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\UARTTransmitter_ins.txCounter[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\SRAMController_ins.sram_tmp[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\UARTTransmitter_ins.txCounter[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\UARTReceiver_ins.inputReg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\UARTReceiver_ins.rxCounter[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\UARTTransmitter_ins.txCounter[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\SRAMController_ins.rx_data_out[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\SRAMController_ins.sram_tmp[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\SRAMController_ins.sram_tmp[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\UARTTransmitter_ins.txCounter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\UARTTransmitter_ins.txCounter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\UARTReceiver_ins.rxCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\UARTReceiver_ins.rxCounter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\UARTReceiver_ins.rxCounter[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\dpu_ins.data_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\UARTReceiver_ins.data[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\UARTTransmitter_ins.txCounter[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\SRAMController_ins.sram_tmp[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\SRAMController_ins.rx_data_out[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\UARTReceiver_ins.data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\UARTReceiver_ins.data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\UARTTransmitter_ins.txCounter[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\UARTReceiver_ins.data[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\SRAMController_ins.sram_tmp[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\UARTReceiver_ins.inputReg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\dpu_ins.data_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_sram_ins_csb0 (.DIODE(\SRAMController_ins.csb_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__X (.DIODE(\SRAMController_ins.csb_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__Q (.DIODE(\SRAMController_ins.data_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A0 (.DIODE(\SRAMController_ins.data_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__A1 (.DIODE(\SRAMController_ins.data_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__A1 (.DIODE(\SRAMController_ins.data_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__Q (.DIODE(\SRAMController_ins.data_tmp[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__A0 (.DIODE(\SRAMController_ins.data_tmp[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A1 (.DIODE(\SRAMController_ins.data_tmp[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1192__A1 (.DIODE(\SRAMController_ins.data_tmp[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__Q (.DIODE(\SRAMController_ins.data_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__A0 (.DIODE(\SRAMController_ins.data_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__A1 (.DIODE(\SRAMController_ins.data_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__A1 (.DIODE(\SRAMController_ins.data_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__Q (.DIODE(\SRAMController_ins.data_tmp[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1546__A0 (.DIODE(\SRAMController_ins.data_tmp[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__A1 (.DIODE(\SRAMController_ins.data_tmp[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__A1 (.DIODE(\SRAMController_ins.data_tmp[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__Q (.DIODE(\SRAMController_ins.data_tmp[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__A0 (.DIODE(\SRAMController_ins.data_tmp[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__A1 (.DIODE(\SRAMController_ins.data_tmp[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__A1 (.DIODE(\SRAMController_ins.data_tmp[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__Q (.DIODE(\SRAMController_ins.data_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__A0 (.DIODE(\SRAMController_ins.data_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1533__A1 (.DIODE(\SRAMController_ins.data_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__A1 (.DIODE(\SRAMController_ins.data_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1770__Q (.DIODE(\SRAMController_ins.data_tmp[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__A0 (.DIODE(\SRAMController_ins.data_tmp[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A1 (.DIODE(\SRAMController_ins.data_tmp[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__A1 (.DIODE(\SRAMController_ins.data_tmp[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1771__Q (.DIODE(\SRAMController_ins.data_tmp[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1554__A0 (.DIODE(\SRAMController_ins.data_tmp[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__A1 (.DIODE(\SRAMController_ins.data_tmp[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__A1 (.DIODE(\SRAMController_ins.data_tmp[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__Q (.DIODE(\SRAMController_ins.data_tmp[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__A0 (.DIODE(\SRAMController_ins.data_tmp[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A1 (.DIODE(\SRAMController_ins.data_tmp[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1199__A1 (.DIODE(\SRAMController_ins.data_tmp[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__Q (.DIODE(\SRAMController_ins.data_tmp[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1558__A0 (.DIODE(\SRAMController_ins.data_tmp[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__A1 (.DIODE(\SRAMController_ins.data_tmp[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1200__A1 (.DIODE(\SRAMController_ins.data_tmp[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1774__Q (.DIODE(\SRAMController_ins.data_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1561__A0 (.DIODE(\SRAMController_ins.data_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__A1 (.DIODE(\SRAMController_ins.data_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1203__A1 (.DIODE(\SRAMController_ins.data_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__Q (.DIODE(\SRAMController_ins.data_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__A0 (.DIODE(\SRAMController_ins.data_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__A1 (.DIODE(\SRAMController_ins.data_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__A1 (.DIODE(\SRAMController_ins.data_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1779__Q (.DIODE(\SRAMController_ins.data_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__A0 (.DIODE(\SRAMController_ins.data_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1554__A1 (.DIODE(\SRAMController_ins.data_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__A1 (.DIODE(\SRAMController_ins.data_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1780__Q (.DIODE(\SRAMController_ins.data_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__A0 (.DIODE(\SRAMController_ins.data_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__A1 (.DIODE(\SRAMController_ins.data_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1209__A1 (.DIODE(\SRAMController_ins.data_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__Q (.DIODE(\SRAMController_ins.data_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__A0 (.DIODE(\SRAMController_ins.data_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1558__A1 (.DIODE(\SRAMController_ins.data_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__A1 (.DIODE(\SRAMController_ins.data_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__Q (.DIODE(\SRAMController_ins.data_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__A0 (.DIODE(\SRAMController_ins.data_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1561__A1 (.DIODE(\SRAMController_ins.data_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1211__A1 (.DIODE(\SRAMController_ins.data_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__Q (.DIODE(\SRAMController_ins.data_tmp[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__A0 (.DIODE(\SRAMController_ins.data_tmp[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__A1 (.DIODE(\SRAMController_ins.data_tmp[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__A1 (.DIODE(\SRAMController_ins.data_tmp[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__Q (.DIODE(\SRAMController_ins.data_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__A0 (.DIODE(\SRAMController_ins.data_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__A1 (.DIODE(\SRAMController_ins.data_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__A1 (.DIODE(\SRAMController_ins.data_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__Q (.DIODE(\SRAMController_ins.data_tmp[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__A0 (.DIODE(\SRAMController_ins.data_tmp[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__A1 (.DIODE(\SRAMController_ins.data_tmp[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__A1 (.DIODE(\SRAMController_ins.data_tmp[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1762__Q (.DIODE(\SRAMController_ins.data_tmp[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A0 (.DIODE(\SRAMController_ins.data_tmp[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__A1 (.DIODE(\SRAMController_ins.data_tmp[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__A1 (.DIODE(\SRAMController_ins.data_tmp[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1763__Q (.DIODE(\SRAMController_ins.data_tmp[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__A0 (.DIODE(\SRAMController_ins.data_tmp[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__A1 (.DIODE(\SRAMController_ins.data_tmp[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__A1 (.DIODE(\SRAMController_ins.data_tmp[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1672__Q (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__A1 (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1436__A1 (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1329__A1 (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__A1 (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__A (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__Q (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__A1 (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1438__A1 (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__A1 (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1305__A1 (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1158__A (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1674__Q (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__A1 (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__A1 (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1333__A1 (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1307__A1 (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__A (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1676__Q (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__A1 (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__A1 (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1337__A1 (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__A2 (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__B (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__B (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1133__A2 (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__A2 (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(\SRAMController_ins.rx_data_out[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1677__Q (.DIODE(\SRAMController_ins.rx_data_out[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__A1 (.DIODE(\SRAMController_ins.rx_data_out[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__A1 (.DIODE(\SRAMController_ins.rx_data_out[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1804__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1805__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1192__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1806__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1808__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1199__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1200__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1795__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1814__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1203__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1815__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1816__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1205__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1209__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1821__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1822__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1211__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1823__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1796__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1824__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1798__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1801__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__Q (.DIODE(\SRAMController_ins.sram_data_from_dpu[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__B2 (.DIODE(\SRAMController_ins.sram_data_from_dpu[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[0]  (.DIODE(\SRAMController_ins.sram_data_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__X (.DIODE(\SRAMController_ins.sram_data_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[1]  (.DIODE(\SRAMController_ins.sram_data_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__X (.DIODE(\SRAMController_ins.sram_data_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[2]  (.DIODE(\SRAMController_ins.sram_data_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__X (.DIODE(\SRAMController_ins.sram_data_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[11]  (.DIODE(\SRAMController_ins.sram_data_out[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__A1 (.DIODE(\SRAMController_ins.sram_data_out[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[13]  (.DIODE(\SRAMController_ins.sram_data_out[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1476__A1 (.DIODE(\SRAMController_ins.sram_data_out[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[16]  (.DIODE(\SRAMController_ins.sram_data_out[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__A1 (.DIODE(\SRAMController_ins.sram_data_out[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[17]  (.DIODE(\SRAMController_ins.sram_data_out[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__A1 (.DIODE(\SRAMController_ins.sram_data_out[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[19]  (.DIODE(\SRAMController_ins.sram_data_out[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1488__A1 (.DIODE(\SRAMController_ins.sram_data_out[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[20]  (.DIODE(\SRAMController_ins.sram_data_out[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__A1 (.DIODE(\SRAMController_ins.sram_data_out[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[21]  (.DIODE(\SRAMController_ins.sram_data_out[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__A1 (.DIODE(\SRAMController_ins.sram_data_out[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[22]  (.DIODE(\SRAMController_ins.sram_data_out[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__A1 (.DIODE(\SRAMController_ins.sram_data_out[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[23]  (.DIODE(\SRAMController_ins.sram_data_out[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A1 (.DIODE(\SRAMController_ins.sram_data_out[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[24]  (.DIODE(\SRAMController_ins.sram_data_out[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1499__A1 (.DIODE(\SRAMController_ins.sram_data_out[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[25]  (.DIODE(\SRAMController_ins.sram_data_out[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__A1 (.DIODE(\SRAMController_ins.sram_data_out[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[26]  (.DIODE(\SRAMController_ins.sram_data_out[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__A1 (.DIODE(\SRAMController_ins.sram_data_out[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[27]  (.DIODE(\SRAMController_ins.sram_data_out[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A1 (.DIODE(\SRAMController_ins.sram_data_out[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[28]  (.DIODE(\SRAMController_ins.sram_data_out[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__A1 (.DIODE(\SRAMController_ins.sram_data_out[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[29]  (.DIODE(\SRAMController_ins.sram_data_out[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__A1 (.DIODE(\SRAMController_ins.sram_data_out[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[2]  (.DIODE(\SRAMController_ins.sram_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__A1 (.DIODE(\SRAMController_ins.sram_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[30]  (.DIODE(\SRAMController_ins.sram_data_out[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A1 (.DIODE(\SRAMController_ins.sram_data_out[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[31]  (.DIODE(\SRAMController_ins.sram_data_out[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A1 (.DIODE(\SRAMController_ins.sram_data_out[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[3]  (.DIODE(\SRAMController_ins.sram_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__A1 (.DIODE(\SRAMController_ins.sram_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[5]  (.DIODE(\SRAMController_ins.sram_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__A1 (.DIODE(\SRAMController_ins.sram_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[6]  (.DIODE(\SRAMController_ins.sram_data_out[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__A1 (.DIODE(\SRAMController_ins.sram_data_out[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[7]  (.DIODE(\SRAMController_ins.sram_data_out[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__A1 (.DIODE(\SRAMController_ins.sram_data_out[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[8]  (.DIODE(\SRAMController_ins.sram_data_out[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__A1 (.DIODE(\SRAMController_ins.sram_data_out[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[9]  (.DIODE(\SRAMController_ins.sram_data_out[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__A1 (.DIODE(\SRAMController_ins.sram_data_out[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1722__Q (.DIODE(\SRAMController_ins.sram_tmp[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__B2 (.DIODE(\SRAMController_ins.sram_tmp[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1449__A0 (.DIODE(\SRAMController_ins.sram_tmp[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__A1 (.DIODE(\SRAMController_ins.sram_tmp[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__Q (.DIODE(\SRAMController_ins.sram_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__B2 (.DIODE(\SRAMController_ins.sram_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__A0 (.DIODE(\SRAMController_ins.sram_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__B2 (.DIODE(\SRAMController_ins.sram_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__Q (.DIODE(\SRAMController_ins.sram_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__B2 (.DIODE(\SRAMController_ins.sram_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1474__A0 (.DIODE(\SRAMController_ins.sram_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__B2 (.DIODE(\SRAMController_ins.sram_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__Q (.DIODE(\SRAMController_ins.sram_tmp[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__B2 (.DIODE(\SRAMController_ins.sram_tmp[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__A0 (.DIODE(\SRAMController_ins.sram_tmp[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__B2 (.DIODE(\SRAMController_ins.sram_tmp[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1737__Q (.DIODE(\SRAMController_ins.sram_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1626__B2 (.DIODE(\SRAMController_ins.sram_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1480__A0 (.DIODE(\SRAMController_ins.sram_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1408__B2 (.DIODE(\SRAMController_ins.sram_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__Q (.DIODE(\SRAMController_ins.sram_tmp[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__B2 (.DIODE(\SRAMController_ins.sram_tmp[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__A0 (.DIODE(\SRAMController_ins.sram_tmp[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__A1 (.DIODE(\SRAMController_ins.sram_tmp[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__Q (.DIODE(\SRAMController_ins.sram_tmp[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__B2 (.DIODE(\SRAMController_ins.sram_tmp[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__A0 (.DIODE(\SRAMController_ins.sram_tmp[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__A1 (.DIODE(\SRAMController_ins.sram_tmp[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__Q (.DIODE(\SRAMController_ins.sram_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__B2 (.DIODE(\SRAMController_ins.sram_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__A0 (.DIODE(\SRAMController_ins.sram_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__A1 (.DIODE(\SRAMController_ins.sram_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__Q (.DIODE(\SRAMController_ins.sram_tmp[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__B2 (.DIODE(\SRAMController_ins.sram_tmp[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__A0 (.DIODE(\SRAMController_ins.sram_tmp[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__A1 (.DIODE(\SRAMController_ins.sram_tmp[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__Q (.DIODE(\SRAMController_ins.sram_tmp[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__B2 (.DIODE(\SRAMController_ins.sram_tmp[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__A0 (.DIODE(\SRAMController_ins.sram_tmp[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__A1 (.DIODE(\SRAMController_ins.sram_tmp[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__Q (.DIODE(\SRAMController_ins.sram_tmp[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__B2 (.DIODE(\SRAMController_ins.sram_tmp[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A0 (.DIODE(\SRAMController_ins.sram_tmp[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__A1 (.DIODE(\SRAMController_ins.sram_tmp[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__Q (.DIODE(\SRAMController_ins.sram_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__B2 (.DIODE(\SRAMController_ins.sram_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1499__A0 (.DIODE(\SRAMController_ins.sram_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__B2 (.DIODE(\SRAMController_ins.sram_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__Q (.DIODE(\SRAMController_ins.sram_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__B2 (.DIODE(\SRAMController_ins.sram_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__A0 (.DIODE(\SRAMController_ins.sram_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__B2 (.DIODE(\SRAMController_ins.sram_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__Q (.DIODE(\SRAMController_ins.sram_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1639__B2 (.DIODE(\SRAMController_ins.sram_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__A0 (.DIODE(\SRAMController_ins.sram_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__B2 (.DIODE(\SRAMController_ins.sram_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__Q (.DIODE(\SRAMController_ins.sram_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__B2 (.DIODE(\SRAMController_ins.sram_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A0 (.DIODE(\SRAMController_ins.sram_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__B2 (.DIODE(\SRAMController_ins.sram_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__Q (.DIODE(\SRAMController_ins.sram_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__B2 (.DIODE(\SRAMController_ins.sram_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__A0 (.DIODE(\SRAMController_ins.sram_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__B2 (.DIODE(\SRAMController_ins.sram_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__Q (.DIODE(\SRAMController_ins.sram_tmp[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__B2 (.DIODE(\SRAMController_ins.sram_tmp[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__A0 (.DIODE(\SRAMController_ins.sram_tmp[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__B2 (.DIODE(\SRAMController_ins.sram_tmp[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__Q (.DIODE(\SRAMController_ins.sram_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__B2 (.DIODE(\SRAMController_ins.sram_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A0 (.DIODE(\SRAMController_ins.sram_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__B2 (.DIODE(\SRAMController_ins.sram_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1753__Q (.DIODE(\SRAMController_ins.sram_tmp[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__B2 (.DIODE(\SRAMController_ins.sram_tmp[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A0 (.DIODE(\SRAMController_ins.sram_tmp[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__B2 (.DIODE(\SRAMController_ins.sram_tmp[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1725__Q (.DIODE(\SRAMController_ins.sram_tmp[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__B2 (.DIODE(\SRAMController_ins.sram_tmp[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__A0 (.DIODE(\SRAMController_ins.sram_tmp[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__A1 (.DIODE(\SRAMController_ins.sram_tmp[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1726__Q (.DIODE(\SRAMController_ins.sram_tmp[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1613__B2 (.DIODE(\SRAMController_ins.sram_tmp[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__A0 (.DIODE(\SRAMController_ins.sram_tmp[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__A1 (.DIODE(\SRAMController_ins.sram_tmp[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__Q (.DIODE(\SRAMController_ins.sram_tmp[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1614__B2 (.DIODE(\SRAMController_ins.sram_tmp[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__A0 (.DIODE(\SRAMController_ins.sram_tmp[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1400__A1 (.DIODE(\SRAMController_ins.sram_tmp[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1728__Q (.DIODE(\SRAMController_ins.sram_tmp[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1615__B2 (.DIODE(\SRAMController_ins.sram_tmp[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__A0 (.DIODE(\SRAMController_ins.sram_tmp[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__A1 (.DIODE(\SRAMController_ins.sram_tmp[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1729__Q (.DIODE(\SRAMController_ins.sram_tmp[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1616__B2 (.DIODE(\SRAMController_ins.sram_tmp[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__A0 (.DIODE(\SRAMController_ins.sram_tmp[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1408__A1 (.DIODE(\SRAMController_ins.sram_tmp[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_sram_ins_web0 (.DIODE(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__X (.DIODE(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__C1 (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__X (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1382__A2 (.DIODE(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__X (.DIODE(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1386__A2 (.DIODE(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__X (.DIODE(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__A2 (.DIODE(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__X (.DIODE(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__A2 (.DIODE(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__X (.DIODE(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__A2 (.DIODE(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__X (.DIODE(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1402__A2 (.DIODE(_0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__X (.DIODE(_0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1406__A2 (.DIODE(_0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__X (.DIODE(_0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1410__A2 (.DIODE(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__X (.DIODE(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__S (.DIODE(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__S (.DIODE(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1490__A (.DIODE(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__A (.DIODE(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1448__A (.DIODE(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__X (.DIODE(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__S (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__S (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__S (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__S (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__S (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__S (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__S (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__S (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__S (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1449__S (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1448__X (.DIODE(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1488__S (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__S (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__S (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__S (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1480__S (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__S (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1476__S (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1474__S (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__S (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__S (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__X (.DIODE(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__S (.DIODE(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__S (.DIODE(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__A (.DIODE(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__A (.DIODE(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__A (.DIODE(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__X (.DIODE(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__S (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__S (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1533__S (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__S (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__S (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__S (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__S (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__S (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__S (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__S (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__X (.DIODE(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1558__S (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__S (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1554__S (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__S (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__S (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__S (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1546__S (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__S (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__S (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__S (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__X (.DIODE(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__S (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__S (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__S (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__S (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__S (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__S (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__S (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__S (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__S (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1561__S (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__X (.DIODE(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__B1 (.DIODE(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__B1 (.DIODE(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__A (.DIODE(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__A (.DIODE(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1608__A (.DIODE(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__Y (.DIODE(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__B1 (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__B1 (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1616__B1 (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1615__B1 (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1614__B1 (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1613__B1 (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__B1 (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__B1 (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__B1 (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__B1 (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1608__X (.DIODE(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__A2 (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__A2 (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__A2 (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1626__A2 (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__A2 (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__A2 (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__A2 (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__A2 (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__A2 (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__A2 (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__X (.DIODE(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__B1 (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__B1 (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__B1 (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__B1 (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1626__B1 (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__B1 (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__B1 (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__B1 (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__B1 (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__B1 (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__X (.DIODE(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__A2 (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__A2 (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1639__A2 (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__A2 (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__A2 (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__A2 (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__A2 (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__A2 (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__A2 (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__A2 (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__X (.DIODE(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__A2 (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__A (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__A (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1325__A (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1284__C1 (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1272__B1 (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__A (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1232__B1 (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__C1 (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__A1 (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__X (.DIODE(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1408__A2 (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__A2 (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1400__A2 (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__A2 (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__A2 (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__A2 (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__A2 (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__A2 (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__A (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__A (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0820__Y (.DIODE(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__B1 (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__B1 (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__B1 (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__B1 (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__B1 (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__B1 (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__B1 (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__B1 (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__A (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__D (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__Y (.DIODE(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__A2 (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__A2 (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0954__A2 (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0949__A2 (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__A2 (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__A2 (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__A2 (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__A2 (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__A2 (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__B2 (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__X (.DIODE(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__B (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__B (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__B (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0912__B (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0911__B (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__B (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0904__B (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__B (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0891__A (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__A (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__X (.DIODE(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__B (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__B (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__B (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__B (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0943__B (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__B (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0929__B (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0920__B (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0895__B (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__A (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__X (.DIODE(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__B (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__B (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__B (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__B (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1011__B (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__B (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__B (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__B1 (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__B1 (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__A (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__X (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__B (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__B (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1062__B (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__B (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__B (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__B (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1006__B1 (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0989__B1 (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__B1 (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__A (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__X (.DIODE(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1107__B (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__B (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__B (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__B (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__B (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__B (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__A2_N (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__B (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__A2 (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__B (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__X (.DIODE(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__B2 (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__B1 (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__B1 (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0954__B1 (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0949__B1 (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__B1 (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__B1 (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__B1 (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__B1 (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__B1 (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__X (.DIODE(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A1 (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__A1 (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1060__A1 (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1048__A1 (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__A1 (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__A1 (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__B1 (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__A1 (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0919__A1 (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0888__B1 (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__X (.DIODE(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__B (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1003__B (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__B (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__B (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0950__B (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0942__B (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__B (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__B (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0893__B (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__B (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0891__X (.DIODE(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__A2 (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__A2 (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__A2 (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__A2 (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__A2 (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__A2 (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__A2 (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0933__A2 (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__A2 (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__A2 (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__X (.DIODE(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__B1 (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__B1 (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__B1 (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__B1 (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__B1 (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__B1 (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__B1 (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0933__B1 (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__B1 (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__B1 (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0901__X (.DIODE(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__A1 (.DIODE(_0533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__A1 (.DIODE(_0533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__A (.DIODE(_0533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0960__B1_N (.DIODE(_0533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__X (.DIODE(_0533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__A2 (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__A2 (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__A2 (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__A2 (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__A2 (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__A2 (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__A2 (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__A2 (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__A2 (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__A2 (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__X (.DIODE(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__B1 (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__B1 (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__B1 (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__B1 (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__B1 (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__B1 (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__B1 (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__B1 (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__B1 (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__B1 (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__X (.DIODE(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1408__B1 (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__B1 (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1400__B1 (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__B1 (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__B1 (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__B1 (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__B1 (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__B1 (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__A2 (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__A0 (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__X (.DIODE(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__A2 (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__A2 (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__A2 (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__A2 (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__A2 (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__A2 (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__A2 (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__A2 (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__A (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__B (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__X (.DIODE(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__A2 (.DIODE(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__A2 (.DIODE(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1201__A (.DIODE(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__A (.DIODE(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__A (.DIODE(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__A2 (.DIODE(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__A2 (.DIODE(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__A2 (.DIODE(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__A2 (.DIODE(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__Y (.DIODE(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__B1 (.DIODE(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__B1 (.DIODE(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__A (.DIODE(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__A (.DIODE(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__A (.DIODE(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__B1 (.DIODE(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__X (.DIODE(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__A2 (.DIODE(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__A2 (.DIODE(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__A2 (.DIODE(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__A (.DIODE(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__A (.DIODE(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__B (.DIODE(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__A (.DIODE(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__X (.DIODE(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__A2 (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1616__A2 (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1615__A2 (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1614__A2 (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1613__A2 (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__A2 (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__A2 (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__A2 (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__A2 (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__A (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__X (.DIODE(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__A2 (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__A2 (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__A2 (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__A2 (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__A2 (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__A2 (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__A2 (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__A2 (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__A2 (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__A2 (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__X (.DIODE(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__B1 (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__B1 (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__B1 (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__B1 (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__B1 (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__B1 (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__B1 (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__B1 (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__B1 (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__B1 (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__X (.DIODE(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_A (.DIODE(\dpu_ins.cur_cmd[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__B1 (.DIODE(\dpu_ins.cur_cmd[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__A (.DIODE(\dpu_ins.cur_cmd[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__Q (.DIODE(\dpu_ins.cur_cmd[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__Q (.DIODE(\dpu_ins.data_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__A1 (.DIODE(\dpu_ins.data_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__B2 (.DIODE(\dpu_ins.data_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__A (.DIODE(\dpu_ins.data_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__A (.DIODE(\dpu_ins.data_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__A1 (.DIODE(\dpu_ins.data_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__Q (.DIODE(\dpu_ins.data_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__A1 (.DIODE(\dpu_ins.data_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__B2 (.DIODE(\dpu_ins.data_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__A (.DIODE(\dpu_ins.data_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__A (.DIODE(\dpu_ins.data_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__A (.DIODE(\dpu_ins.data_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__A1 (.DIODE(\dpu_ins.data_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__D (.DIODE(\dpu_ins.data_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__X (.DIODE(\dpu_ins.data_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_A (.DIODE(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_A (.DIODE(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_A (.DIODE(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1814__RESET_B (.DIODE(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__A2 (.DIODE(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire3_X (.DIODE(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__A2 (.DIODE(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__A2 (.DIODE(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__B (.DIODE(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout10_X (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__A (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A_N (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__A0 (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__A2_N (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0883__A (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0899__B1 (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__A (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__B1 (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__B1 (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_X (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__A (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__B1 (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1042__A (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1065__B1 (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1080__B1 (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__B1 (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__B1 (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__A (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout10_A (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout11_A (.DIODE(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_X (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__RESET_B (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__RESET_B (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__RESET_B (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_A (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__RESET_B (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__RESET_B (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1780__RESET_B (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_X (.DIODE(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__RESET_B (.DIODE(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__RESET_B (.DIODE(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1760__RESET_B (.DIODE(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__RESET_B (.DIODE(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__RESET_B (.DIODE(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__RESET_B (.DIODE(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_A (.DIODE(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_X (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1721__RESET_B (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1720__RESET_B (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1432__A (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__A (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1316__A (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__A (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1222__A (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0842__A1 (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__A (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout29_X (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1415__A (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__C1 (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__C1 (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_A (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__RESET_B (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1714__RESET_B (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__RESET_B (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout33_X (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout32_A (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__RESET_B (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__RESET_B (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__RESET_B (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__RESET_B (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__RESET_B (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__RESET_B (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1726__RESET_B (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__RESET_B (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1722__RESET_B (.DIODE(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_X (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_A (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__RESET_B (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__RESET_B (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout33_A (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_A (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout30_A (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__RESET_B (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_X (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__RESET_B (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__RESET_B (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__RESET_B (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__RESET_B (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1753__RESET_B (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__RESET_B (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout35_A (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__RESET_B (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__RESET_B (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1843__RESET_B (.DIODE(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_X (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__RESET_B (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__RESET_B (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__RESET_B (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__RESET_B (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__RESET_B (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__RESET_B (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__RESET_B (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1737__RESET_B (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__RESET_B (.DIODE(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_X (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__RESET_B (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__RESET_B (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__RESET_B (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__RESET_B (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__RESET_B (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__RESET_B (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__RESET_B (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1774__RESET_B (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__RESET_B (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__RESET_B (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_X (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__RESET_B (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__RESET_B (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1824__RESET_B (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1823__RESET_B (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1822__RESET_B (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1821__RESET_B (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__RESET_B (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_A (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__RESET_B (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__RESET_B (.DIODE(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_X (.DIODE(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__RESET_B (.DIODE(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__RESET_B (.DIODE(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__RESET_B (.DIODE(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_A (.DIODE(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__RESET_B (.DIODE(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__RESET_B (.DIODE(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__RESET_B (.DIODE(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__RESET_B (.DIODE(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1694__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1701__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1706__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1689__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1686__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1707__CLK (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_X (.DIODE(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload6_A (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1837__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1806__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1805__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1804__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1731__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1801__CLK (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_X (.DIODE(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload13_A (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1822__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1821__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1824__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1852__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1851__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1816__CLK (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_X (.DIODE(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload16_A (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__CLK (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__CLK (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__CLK (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__CLK (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__CLK (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1774__CLK (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__CLK (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__CLK (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__CLK (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_X (.DIODE(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload17_A (.DIODE(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__CLK (.DIODE(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__CLK (.DIODE(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1726__CLK (.DIODE(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__CLK (.DIODE(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__CLK (.DIODE(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__CLK (.DIODE(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1737__CLK (.DIODE(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__CLK (.DIODE(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_X (.DIODE(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_clk_X (.DIODE(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload0_A (.DIODE(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_clk_X (.DIODE(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\SRAMController_ins.sram_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\SRAMController_ins.sram_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\SRAMController_ins.sram_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\SRAMController_ins.sram_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\SRAMController_ins.sram_data_from_dpu[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\SRAMController_ins.sram_data_out[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\SRAMController_ins.sram_data_out[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_234 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_454 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_487 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_595 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_619 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_647 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_659 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_667 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_716 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_735 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_742 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_752 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_767 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_783 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_798 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_828 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_883 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_901 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_907 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_919 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_957 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_965 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1006 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_507 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_524 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_599 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_716 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_736 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_766 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1003 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1034 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1046 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1058 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_451 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_472 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_488 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_570 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_621 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_639 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_647 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_650 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_660 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_688 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_714 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_729 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_741 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_777 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_859 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_884 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_912 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_920 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_959 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1034 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1018 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1030 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1066 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1030 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1038 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1018 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1030 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1066 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1025 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1018 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1030 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1066 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1018 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1030 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1038 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1027 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1039 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1051 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1031 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1039 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1041 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1053 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1065 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1018 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1030 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1038 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1031 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1039 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1031 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1043 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1055 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1067 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1031 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1043 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1055 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1067 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1031 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1039 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_140 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_152 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_151 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_99 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_79 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_91 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_172 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_49 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_112 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_124 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_92 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_144 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_87 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_42 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_54 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_66 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_101 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_172 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_173 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_110 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_33 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_100 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_112 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_55 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_67 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_152 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1022 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1034 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_119 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_131 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_369 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_434 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_449 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_461 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_499 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_514 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_561 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_573 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_645 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_657 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_673 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_723 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_759 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_787 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_815 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_821 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_841 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_853 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_978 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_981 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_993 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_472 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_661 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_766 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_778 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_795 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_803 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_849 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_879 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_885 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_890 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_901 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_938 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_950 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_961 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_984 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_996 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1033 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1045 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_205 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_431 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_479 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_598 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_621 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_649 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_652 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_722 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_765 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_807 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_859 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_900 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_912 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_927 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_935 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1006 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1018 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1030 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1061 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1073 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_42 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_339 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_403 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_457 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_492 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_516 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_526 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_539 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_626 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_694 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_719 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_731 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_758 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_764 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_779 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_793 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_805 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_826 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_831 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_837 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_863 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_934 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_943 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_965 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_972 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_976 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_983 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_994 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1006 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1033 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1045 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_199 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_350 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_459 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_467 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_481 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_493 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_505 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_517 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_537 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_582 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_610 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_619 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_623 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_649 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_696 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_718 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_739 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_754 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_771 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_778 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_789 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_835 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_881 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_894 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_906 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_914 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_933 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_946 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_954 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_996 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1008 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1020 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1032 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1061 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1073 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_484 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_535 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_588 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_666 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_694 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_704 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_723 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_731 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_743 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_751 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_764 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_800 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_812 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_818 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_852 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_860 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_863 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_881 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_885 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_889 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_892 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_911 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_915 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_946 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_967 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_996 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1033 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1045 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_146 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_708 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_741 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_751 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_773 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_792 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_801 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_809 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_849 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_858 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_862 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_952 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_981 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_993 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1005 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1017 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1029 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1061 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1073 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_155 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_227 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_267 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_366 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_482 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_520 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_546 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_623 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_675 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_696 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_713 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_756 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_760 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_789 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_802 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_891 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_912 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_924 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_930 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_950 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_978 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_990 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1002 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1033 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1045 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_154 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_203 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_225 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_237 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_311 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_323 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_339 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_351 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_393 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_405 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_460 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_472 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_489 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_499 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_505 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_517 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_549 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_571 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_617 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_647 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_659 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_668 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_682 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_694 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_713 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_729 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_741 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_753 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_769 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_777 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_781 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_785 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_797 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_809 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_813 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_825 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_837 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_843 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_847 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_859 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_864 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_879 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_891 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_897 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_909 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_925 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_937 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_953 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_965 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_981 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_993 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 assign uio_oe[0] = net47;
 assign uio_oe[1] = net48;
 assign uio_oe[2] = net49;
 assign uio_oe[3] = net50;
 assign uio_oe[4] = net67;
 assign uio_oe[5] = net51;
 assign uio_oe[6] = net52;
 assign uio_oe[7] = net53;
 assign uio_out[0] = net54;
 assign uio_out[1] = net55;
 assign uio_out[2] = net56;
 assign uio_out[3] = net57;
 assign uio_out[5] = net58;
 assign uio_out[6] = net59;
 assign uio_out[7] = net60;
 assign uo_out[1] = net61;
 assign uo_out[2] = net62;
 assign uo_out[3] = net63;
 assign uo_out[4] = net64;
 assign uo_out[5] = net65;
endmodule
