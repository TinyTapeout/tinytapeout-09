MACRO tt_um_urish_charge_pump
  CLASS BLOCK ;
  FOREIGN tt_um_urish_charge_pump ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.804199 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 25.734600 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 126.560 5.000 128.060 220.760 ;
    END
  END VAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 33.360 5.000 34.860 220.760 ;
    END
  END VGND
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.360 5.000 31.860 220.760 ;
    END
  END VDPWR
  OBS
      LAYER pwell ;
        RECT 135.800 220.490 138.580 224.070 ;
        RECT 135.800 216.350 138.580 219.930 ;
      LAYER nwell ;
        RECT 138.830 215.600 141.910 224.210 ;
      LAYER pwell ;
        RECT 90.260 212.420 95.040 213.320 ;
        RECT 90.260 209.440 91.160 212.420 ;
      LAYER nwell ;
        RECT 91.160 209.440 94.140 212.420 ;
      LAYER pwell ;
        RECT 94.140 209.440 95.040 212.420 ;
        RECT 90.260 208.540 95.040 209.440 ;
        RECT 90.300 184.310 95.080 185.210 ;
        RECT 90.300 181.330 91.200 184.310 ;
      LAYER nwell ;
        RECT 91.200 181.330 94.180 184.310 ;
      LAYER pwell ;
        RECT 94.180 181.330 95.080 184.310 ;
        RECT 90.300 180.430 95.080 181.330 ;
        RECT 90.270 157.270 95.050 158.170 ;
        RECT 90.270 154.290 91.170 157.270 ;
      LAYER nwell ;
        RECT 91.170 154.290 94.150 157.270 ;
      LAYER pwell ;
        RECT 94.150 154.290 95.050 157.270 ;
        RECT 90.270 153.390 95.050 154.290 ;
        RECT 90.270 140.850 95.050 141.750 ;
        RECT 90.270 137.870 91.170 140.850 ;
      LAYER nwell ;
        RECT 91.170 137.870 94.150 140.850 ;
      LAYER pwell ;
        RECT 94.150 137.870 95.050 140.850 ;
        RECT 90.270 136.970 95.050 137.870 ;
      LAYER nwell ;
        RECT 100.360 18.050 142.940 21.440 ;
        RECT 100.360 12.480 142.940 15.870 ;
        RECT 100.360 7.000 142.940 10.390 ;
      LAYER li1 ;
        RECT 136.040 223.660 138.340 223.830 ;
        RECT 136.040 220.900 136.210 223.660 ;
        RECT 136.940 222.970 137.440 223.140 ;
        RECT 136.710 221.760 136.880 222.800 ;
        RECT 137.500 221.760 137.670 222.800 ;
        RECT 136.940 221.420 137.440 221.590 ;
        RECT 138.170 220.900 138.340 223.660 ;
        RECT 136.040 220.730 138.340 220.900 ;
        RECT 139.220 223.650 141.520 223.820 ;
        RECT 139.220 220.300 139.390 223.650 ;
        RECT 141.350 223.340 141.520 223.650 ;
        RECT 140.120 222.960 140.620 223.130 ;
        RECT 139.890 221.205 140.060 222.745 ;
        RECT 140.680 221.205 140.850 222.745 ;
        RECT 140.120 220.820 140.620 220.990 ;
        RECT 141.340 220.600 141.520 223.340 ;
        RECT 141.350 220.300 141.520 220.600 ;
        RECT 139.220 220.130 141.520 220.300 ;
        RECT 136.040 219.520 138.340 219.690 ;
        RECT 136.040 216.760 136.210 219.520 ;
        RECT 136.940 218.830 137.440 219.000 ;
        RECT 136.710 217.620 136.880 218.660 ;
        RECT 137.500 217.620 137.670 218.660 ;
        RECT 136.940 217.280 137.440 217.450 ;
        RECT 138.170 216.760 138.340 219.520 ;
        RECT 136.040 216.590 138.340 216.760 ;
        RECT 139.220 219.510 141.520 219.680 ;
        RECT 139.220 216.160 139.390 219.510 ;
        RECT 141.350 219.220 141.520 219.510 ;
        RECT 140.120 218.820 140.620 218.990 ;
        RECT 139.890 217.065 140.060 218.605 ;
        RECT 140.680 217.065 140.850 218.605 ;
        RECT 140.120 216.680 140.620 216.850 ;
        RECT 141.340 216.480 141.520 219.220 ;
        RECT 141.350 216.160 141.520 216.480 ;
        RECT 139.220 215.990 141.520 216.160 ;
        RECT 90.500 213.020 94.800 213.080 ;
        RECT 90.280 212.910 94.800 213.020 ;
        RECT 90.280 208.950 90.970 212.910 ;
        RECT 91.550 211.860 93.750 212.030 ;
        RECT 91.550 210.000 91.720 211.860 ;
        RECT 92.130 210.490 93.170 211.370 ;
        RECT 93.580 211.360 93.750 211.860 ;
        RECT 93.540 210.620 93.780 211.360 ;
        RECT 93.580 210.000 93.750 210.620 ;
        RECT 91.550 209.830 93.750 210.000 ;
        RECT 94.630 208.950 94.800 212.910 ;
        RECT 90.280 208.900 94.800 208.950 ;
        RECT 90.500 208.780 94.800 208.900 ;
        RECT 90.540 184.900 94.840 184.970 ;
        RECT 90.280 184.800 94.840 184.900 ;
        RECT 90.280 180.840 90.970 184.800 ;
        RECT 91.590 183.750 93.790 183.920 ;
        RECT 91.590 181.890 91.760 183.750 ;
        RECT 93.620 183.280 93.790 183.750 ;
        RECT 92.170 182.380 93.210 183.260 ;
        RECT 93.570 182.420 93.880 183.280 ;
        RECT 93.620 181.890 93.790 182.420 ;
        RECT 91.590 181.720 93.790 181.890 ;
        RECT 94.670 180.840 94.840 184.800 ;
        RECT 90.280 180.780 94.840 180.840 ;
        RECT 90.540 180.670 94.840 180.780 ;
        RECT 90.510 157.840 94.810 157.930 ;
        RECT 90.300 157.760 94.810 157.840 ;
        RECT 90.300 153.800 90.990 157.760 ;
        RECT 91.560 156.710 93.760 156.880 ;
        RECT 91.560 154.850 91.730 156.710 ;
        RECT 93.590 156.300 93.760 156.710 ;
        RECT 92.140 155.340 93.180 156.220 ;
        RECT 93.580 155.410 93.780 156.300 ;
        RECT 93.590 154.850 93.760 155.410 ;
        RECT 91.560 154.680 93.760 154.850 ;
        RECT 94.640 153.800 94.810 157.760 ;
        RECT 90.300 153.720 94.810 153.800 ;
        RECT 90.510 153.630 94.810 153.720 ;
        RECT 90.940 141.510 94.400 141.710 ;
        RECT 90.510 141.340 94.810 141.510 ;
        RECT 90.510 137.380 90.680 141.340 ;
        RECT 90.940 141.240 94.400 141.340 ;
        RECT 91.480 140.290 93.760 140.460 ;
        RECT 91.480 138.430 91.780 140.290 ;
        RECT 92.140 138.920 93.180 139.800 ;
        RECT 93.590 138.430 93.760 140.290 ;
        RECT 91.480 138.320 93.760 138.430 ;
        RECT 91.560 138.260 93.760 138.320 ;
        RECT 94.640 137.380 94.810 141.340 ;
        RECT 90.510 137.210 94.810 137.380 ;
        RECT 140.160 21.050 142.130 21.070 ;
        RECT 100.750 20.880 142.550 21.050 ;
        RECT 100.750 18.610 100.920 20.880 ;
        RECT 140.160 20.850 142.130 20.880 ;
        RECT 101.650 20.190 141.650 20.360 ;
        RECT 101.420 19.515 101.590 19.975 ;
        RECT 141.710 19.515 141.880 19.975 ;
        RECT 101.650 19.130 141.650 19.300 ;
        RECT 142.380 18.610 142.550 20.880 ;
        RECT 100.750 18.440 142.550 18.610 ;
        RECT 101.250 15.480 102.650 15.560 ;
        RECT 100.750 15.310 142.550 15.480 ;
        RECT 100.750 13.040 100.920 15.310 ;
        RECT 101.250 15.230 102.650 15.310 ;
        RECT 101.650 14.620 141.650 14.790 ;
        RECT 101.420 13.945 101.590 14.405 ;
        RECT 141.710 13.945 141.880 14.405 ;
        RECT 101.650 13.560 141.650 13.730 ;
        RECT 142.380 13.040 142.550 15.310 ;
        RECT 100.750 12.870 142.550 13.040 ;
        RECT 100.750 9.830 142.550 10.000 ;
        RECT 100.750 7.560 100.920 9.830 ;
        RECT 101.650 9.140 141.650 9.310 ;
        RECT 101.420 8.465 101.590 8.925 ;
        RECT 141.710 8.465 141.880 8.925 ;
        RECT 101.650 8.080 141.650 8.250 ;
        RECT 142.380 7.560 142.550 9.830 ;
        RECT 100.750 7.390 142.550 7.560 ;
      LAYER met1 ;
        RECT 136.960 223.130 137.420 223.170 ;
        RECT 138.110 223.130 138.510 223.180 ;
        RECT 140.140 223.130 140.600 223.160 ;
        RECT 136.960 222.960 140.600 223.130 ;
        RECT 136.960 222.940 137.420 222.960 ;
        RECT 138.110 222.920 138.510 222.960 ;
        RECT 140.140 222.930 140.600 222.960 ;
        RECT 136.490 222.780 136.790 222.810 ;
        RECT 135.970 221.700 136.280 221.800 ;
        RECT 136.490 221.780 136.910 222.780 ;
        RECT 137.470 222.370 137.700 222.780 ;
        RECT 140.770 222.725 141.580 223.560 ;
        RECT 139.860 222.370 140.090 222.725 ;
        RECT 137.470 222.070 140.090 222.370 ;
        RECT 137.470 221.780 137.700 222.070 ;
        RECT 136.490 221.700 136.790 221.780 ;
        RECT 130.110 221.400 136.790 221.700 ;
        RECT 135.970 221.250 136.280 221.400 ;
        RECT 136.960 221.390 137.420 221.620 ;
        RECT 138.160 219.900 138.460 222.070 ;
        RECT 139.860 221.225 140.090 222.070 ;
        RECT 140.650 221.225 141.580 222.725 ;
        RECT 140.140 220.790 140.600 221.020 ;
        RECT 138.110 219.600 138.510 219.900 ;
        RECT 138.160 219.160 138.460 219.600 ;
        RECT 136.940 218.860 140.620 219.160 ;
        RECT 136.960 218.800 137.420 218.860 ;
        RECT 140.140 218.790 140.600 218.860 ;
        RECT 136.010 218.400 136.240 218.460 ;
        RECT 136.680 218.400 136.910 218.640 ;
        RECT 130.110 218.100 136.910 218.400 ;
        RECT 136.010 218.040 136.240 218.100 ;
        RECT 136.680 217.640 136.910 218.100 ;
        RECT 137.470 218.000 137.700 218.640 ;
        RECT 140.770 218.585 141.580 221.225 ;
        RECT 139.860 218.000 140.090 218.585 ;
        RECT 137.470 217.700 140.090 218.000 ;
        RECT 137.470 217.640 138.060 217.700 ;
        RECT 137.520 217.620 138.060 217.640 ;
        RECT 136.960 217.250 137.420 217.480 ;
        RECT 137.760 215.700 138.060 217.620 ;
        RECT 139.860 217.085 140.090 217.700 ;
        RECT 140.650 217.085 141.580 218.585 ;
        RECT 140.140 216.650 140.600 216.880 ;
        RECT 140.770 216.420 141.580 217.085 ;
        RECT 137.610 214.800 138.310 215.700 ;
        RECT 90.250 213.020 91.000 213.080 ;
        RECT 90.230 208.900 91.020 213.020 ;
        RECT 92.150 210.460 93.150 211.400 ;
        RECT 93.510 211.370 93.810 211.420 ;
        RECT 95.190 211.370 96.910 211.500 ;
        RECT 93.510 210.600 96.910 211.370 ;
        RECT 93.510 210.560 93.810 210.600 ;
        RECT 90.250 208.840 91.000 208.900 ;
        RECT 90.250 184.900 91.000 184.960 ;
        RECT 90.230 180.780 91.020 184.900 ;
        RECT 93.540 183.300 93.910 183.340 ;
        RECT 92.190 183.280 93.190 183.290 ;
        RECT 92.190 182.380 93.200 183.280 ;
        RECT 93.540 182.400 96.910 183.300 ;
        RECT 92.190 182.350 93.190 182.380 ;
        RECT 93.540 182.360 93.910 182.400 ;
        RECT 90.250 180.720 91.000 180.780 ;
        RECT 90.270 157.840 91.020 157.900 ;
        RECT 90.250 153.720 91.040 157.840 ;
        RECT 93.550 156.300 93.810 156.360 ;
        RECT 92.160 155.310 93.160 156.250 ;
        RECT 93.550 155.400 96.930 156.300 ;
        RECT 93.550 155.350 93.810 155.400 ;
        RECT 90.270 153.660 91.020 153.720 ;
        RECT 90.080 141.770 95.000 141.780 ;
        RECT 90.070 141.130 95.000 141.770 ;
        RECT 90.080 141.060 95.000 141.130 ;
        RECT 81.260 140.730 85.460 141.000 ;
        RECT 81.260 140.700 91.840 140.730 ;
        RECT 81.210 139.500 91.840 140.700 ;
        RECT 81.260 138.300 91.840 139.500 ;
        RECT 92.150 138.930 93.160 139.830 ;
        RECT 92.160 138.890 93.160 138.930 ;
        RECT 81.210 138.050 91.840 138.300 ;
        RECT 81.210 137.100 85.460 138.050 ;
        RECT 81.260 135.900 85.460 137.100 ;
        RECT 81.210 134.700 85.460 135.900 ;
        RECT 81.260 134.400 85.460 134.700 ;
        RECT 141.570 21.100 142.630 21.350 ;
        RECT 140.100 20.820 142.640 21.100 ;
        RECT 141.570 20.760 142.640 20.820 ;
        RECT 101.210 20.160 141.630 20.390 ;
        RECT 101.210 19.330 102.650 20.160 ;
        RECT 141.780 19.955 142.640 20.760 ;
        RECT 141.680 19.535 142.640 19.955 ;
        RECT 101.210 19.100 141.630 19.330 ;
        RECT 141.780 19.210 142.640 19.535 ;
        RECT 101.210 15.590 102.650 19.100 ;
        RECT 101.190 15.200 102.710 15.590 ;
        RECT 101.210 15.050 102.650 15.200 ;
        RECT 101.210 14.385 101.460 15.050 ;
        RECT 101.670 14.590 141.630 14.820 ;
        RECT 141.810 14.385 142.010 14.510 ;
        RECT 101.210 13.965 101.620 14.385 ;
        RECT 141.680 13.965 142.010 14.385 ;
        RECT 101.210 13.870 101.460 13.965 ;
        RECT 141.810 13.760 142.010 13.965 ;
        RECT 101.670 13.530 142.010 13.760 ;
        RECT 141.810 11.960 142.010 13.530 ;
        RECT 141.660 11.230 142.100 11.960 ;
        RECT 141.810 10.030 142.010 11.230 ;
        RECT 141.750 9.800 142.070 10.030 ;
        RECT 101.670 9.320 141.630 9.340 ;
        RECT 101.330 9.110 141.630 9.320 ;
        RECT 101.330 8.280 101.840 9.110 ;
        RECT 141.810 8.905 142.010 9.800 ;
        RECT 141.680 8.485 142.010 8.905 ;
        RECT 101.330 8.050 141.630 8.280 ;
        RECT 101.330 5.660 101.840 8.050 ;
        RECT 141.810 7.590 142.010 8.485 ;
        RECT 141.750 7.360 142.070 7.590 ;
        RECT 101.330 5.160 101.850 5.660 ;
        RECT 101.330 5.100 101.840 5.160 ;
      LAYER met2 ;
        RECT 128.110 224.660 128.610 225.260 ;
        RECT 128.210 224.410 128.510 224.660 ;
        RECT 128.210 224.110 138.460 224.410 ;
        RECT 138.160 222.870 138.460 224.110 ;
        RECT 130.160 221.350 131.060 221.750 ;
        RECT 123.860 219.900 124.460 219.950 ;
        RECT 138.160 219.900 138.460 219.950 ;
        RECT 123.860 219.300 138.560 219.900 ;
        RECT 123.860 219.250 124.460 219.300 ;
        RECT 130.160 218.050 131.060 218.450 ;
        RECT 13.960 217.710 18.160 217.990 ;
        RECT 13.400 217.430 18.160 217.710 ;
        RECT 12.840 217.150 18.160 217.430 ;
        RECT 12.280 216.870 18.160 217.150 ;
        RECT 12.000 216.590 18.160 216.870 ;
        RECT 11.720 216.310 18.160 216.590 ;
        RECT 20.960 216.310 23.760 217.430 ;
        RECT 11.440 216.030 18.160 216.310 ;
        RECT 11.160 215.470 18.160 216.030 ;
        RECT 10.880 214.910 18.160 215.470 ;
        RECT 10.600 214.630 18.160 214.910 ;
        RECT 21.240 214.630 24.040 216.310 ;
        RECT 10.600 214.350 14.800 214.630 ;
        RECT 10.320 214.070 13.960 214.350 ;
        RECT 10.320 213.790 13.680 214.070 ;
        RECT 10.320 213.510 13.400 213.790 ;
        RECT 10.320 212.950 13.120 213.510 ;
        RECT 10.320 211.550 12.840 212.950 ;
        RECT 10.320 210.710 13.120 211.550 ;
        RECT 10.320 210.430 13.400 210.710 ;
        RECT 10.600 210.150 13.680 210.430 ;
        RECT 10.600 209.870 13.960 210.150 ;
        RECT 10.600 209.590 14.520 209.870 ;
        RECT 15.640 209.590 18.160 214.630 ;
        RECT 21.520 212.110 24.320 214.630 ;
        RECT 21.240 211.270 24.320 212.110 ;
        RECT 20.960 210.710 24.320 211.270 ;
        RECT 20.680 210.430 24.040 210.710 ;
        RECT 20.400 210.150 24.040 210.430 ;
        RECT 20.120 209.870 24.040 210.150 ;
        RECT 19.560 209.590 24.040 209.870 ;
        RECT 10.880 209.310 18.160 209.590 ;
        RECT 19.000 209.310 23.760 209.590 ;
        RECT 10.880 209.030 23.760 209.310 ;
        RECT 11.160 208.470 23.480 209.030 ;
        RECT 90.280 208.850 90.970 213.070 ;
        RECT 92.210 210.470 93.060 211.420 ;
        RECT 11.440 208.190 23.200 208.470 ;
        RECT 11.720 207.910 22.920 208.190 ;
        RECT 12.000 207.630 22.640 207.910 ;
        RECT 12.280 207.350 22.640 207.630 ;
        RECT 12.560 207.070 22.080 207.350 ;
        RECT 13.120 206.790 21.800 207.070 ;
        RECT 13.680 206.510 21.240 206.790 ;
        RECT 14.240 206.230 20.680 206.510 ;
        RECT 15.360 205.950 19.840 206.230 ;
        RECT 10.600 202.030 13.120 203.990 ;
        RECT 24.320 203.710 25.440 203.990 ;
        RECT 23.480 203.430 26.560 203.710 ;
        RECT 22.920 203.150 27.120 203.430 ;
        RECT 22.640 202.870 27.400 203.150 ;
        RECT 22.360 202.590 27.680 202.870 ;
        RECT 13.960 202.310 15.920 202.590 ;
        RECT 22.080 202.310 27.960 202.590 ;
        RECT 13.400 202.030 17.040 202.310 ;
        RECT 22.080 202.030 28.240 202.310 ;
        RECT 10.600 201.750 17.600 202.030 ;
        RECT 21.800 201.750 28.240 202.030 ;
        RECT 10.600 201.470 17.880 201.750 ;
        RECT 21.800 201.470 28.520 201.750 ;
        RECT 10.600 201.190 18.160 201.470 ;
        RECT 10.600 200.910 18.440 201.190 ;
        RECT 10.600 200.350 18.720 200.910 ;
        RECT 21.520 200.630 28.800 201.470 ;
        RECT 21.520 200.350 29.080 200.630 ;
        RECT 10.600 199.790 19.000 200.350 ;
        RECT 21.240 200.070 24.880 200.350 ;
        RECT 25.720 200.070 29.080 200.350 ;
        RECT 10.600 199.230 19.280 199.790 ;
        RECT 10.320 198.950 13.960 199.230 ;
        RECT 15.920 198.950 19.280 199.230 ;
        RECT 21.240 199.510 24.320 200.070 ;
        RECT 26.000 199.790 29.080 200.070 ;
        RECT 26.280 199.510 29.360 199.790 ;
        RECT 10.320 198.670 13.400 198.950 ;
        RECT 16.480 198.670 19.560 198.950 ;
        RECT 10.320 198.110 13.120 198.670 ;
        RECT 16.760 198.110 19.560 198.670 ;
        RECT 10.320 196.150 12.840 198.110 ;
        RECT 17.040 196.150 19.560 198.110 ;
        RECT 10.320 195.590 13.120 196.150 ;
        RECT 16.760 195.590 19.560 196.150 ;
        RECT 21.240 198.110 24.040 199.510 ;
        RECT 26.560 198.950 29.360 199.510 ;
        RECT 21.240 195.590 23.760 198.110 ;
        RECT 26.840 197.550 29.360 198.950 ;
        RECT 27.120 196.710 29.360 197.550 ;
        RECT 10.320 195.310 13.400 195.590 ;
        RECT 16.480 195.310 19.280 195.590 ;
        RECT 10.600 195.030 13.960 195.310 ;
        RECT 15.920 195.030 19.280 195.310 ;
        RECT 20.960 195.310 24.040 195.590 ;
        RECT 26.840 195.310 29.360 196.710 ;
        RECT 20.960 195.030 24.320 195.310 ;
        RECT 10.600 194.750 19.560 195.030 ;
        RECT 20.680 194.750 24.320 195.030 ;
        RECT 26.560 194.750 29.360 195.310 ;
        RECT 10.600 194.470 19.840 194.750 ;
        RECT 20.120 194.470 24.880 194.750 ;
        RECT 26.280 194.470 29.360 194.750 ;
        RECT 10.880 194.190 29.360 194.470 ;
        RECT 10.880 193.910 29.080 194.190 ;
        RECT 11.160 193.350 29.080 193.910 ;
        RECT 11.440 193.070 28.800 193.350 ;
        RECT 11.720 192.790 28.800 193.070 ;
        RECT 12.000 192.510 28.800 192.790 ;
        RECT 12.560 192.230 17.320 192.510 ;
        RECT 18.440 192.230 22.920 192.510 ;
        RECT 23.200 192.230 28.520 192.510 ;
        RECT 12.840 191.950 17.040 192.230 ;
        RECT 18.720 191.950 22.640 192.230 ;
        RECT 13.960 191.670 16.200 191.950 ;
        RECT 19.280 191.670 22.080 191.950 ;
        RECT 23.480 191.670 28.240 192.230 ;
        RECT 20.120 191.390 21.520 191.670 ;
        RECT 24.040 191.390 27.960 191.670 ;
        RECT 24.320 191.110 27.400 191.390 ;
        RECT 24.880 190.830 26.840 191.110 ;
        RECT 13.400 188.030 24.040 188.310 ;
        RECT 12.560 187.750 24.040 188.030 ;
        RECT 12.000 187.470 24.040 187.750 ;
        RECT 11.720 187.190 24.040 187.470 ;
        RECT 11.440 186.910 24.040 187.190 ;
        RECT 11.160 186.630 24.040 186.910 ;
        RECT 95.960 186.720 96.860 211.550 ;
        RECT 10.880 186.070 24.040 186.630 ;
        RECT 10.600 185.230 24.040 186.070 ;
        RECT 92.170 185.820 96.860 186.720 ;
        RECT 10.600 184.950 22.640 185.230 ;
        RECT 10.320 184.670 14.520 184.950 ;
        RECT 10.320 184.390 13.680 184.670 ;
        RECT 10.320 183.830 13.400 184.390 ;
        RECT 10.320 183.270 13.120 183.830 ;
        RECT 10.320 181.030 12.840 183.270 ;
        RECT 15.640 181.870 18.160 184.950 ;
        RECT 19.840 184.670 22.920 184.950 ;
        RECT 20.120 184.390 23.200 184.670 ;
        RECT 20.400 183.830 23.480 184.390 ;
        RECT 20.680 183.550 23.760 183.830 ;
        RECT 20.960 183.270 23.760 183.550 ;
        RECT 21.240 182.710 24.040 183.270 ;
        RECT 21.520 182.150 24.040 182.710 ;
        RECT 15.640 181.310 18.440 181.870 ;
        RECT 21.520 181.310 24.320 182.150 ;
        RECT 15.640 181.030 18.720 181.310 ;
        RECT 10.320 179.910 13.120 181.030 ;
        RECT 15.920 180.750 18.720 181.030 ;
        RECT 21.240 180.750 24.320 181.310 ;
        RECT 15.920 180.470 19.000 180.750 ;
        RECT 20.960 180.470 24.320 180.750 ;
        RECT 90.280 180.730 90.970 184.950 ;
        RECT 92.170 183.330 93.070 185.820 ;
        RECT 92.170 182.370 93.150 183.330 ;
        RECT 92.250 182.330 93.150 182.370 ;
        RECT 15.920 180.190 19.560 180.470 ;
        RECT 20.400 180.190 24.320 180.470 ;
        RECT 15.920 179.910 24.320 180.190 ;
        RECT 10.600 179.630 13.120 179.910 ;
        RECT 16.200 179.630 24.320 179.910 ;
        RECT 10.600 178.790 13.400 179.630 ;
        RECT 16.200 179.070 24.040 179.630 ;
        RECT 16.480 178.790 24.040 179.070 ;
        RECT 10.880 178.230 13.680 178.790 ;
        RECT 16.480 178.510 23.760 178.790 ;
        RECT 16.760 178.230 23.760 178.510 ;
        RECT 10.880 177.950 13.960 178.230 ;
        RECT 17.040 177.950 23.480 178.230 ;
        RECT 11.160 177.670 13.960 177.950 ;
        RECT 17.320 177.670 23.200 177.950 ;
        RECT 17.600 177.390 22.920 177.670 ;
        RECT 17.880 177.110 22.640 177.390 ;
        RECT 18.440 176.830 22.080 177.110 ;
        RECT 19.280 176.550 20.680 176.830 ;
        RECT 10.600 168.430 13.120 173.470 ;
        RECT 20.960 173.190 24.040 173.470 ;
        RECT 21.240 171.790 24.040 173.190 ;
        RECT 21.520 169.830 24.320 171.790 ;
        RECT 21.240 169.270 24.320 169.830 ;
        RECT 20.960 168.990 24.320 169.270 ;
        RECT 20.680 168.710 24.320 168.990 ;
        RECT 20.120 168.430 24.320 168.710 ;
        RECT 6.400 167.310 24.040 168.430 ;
        RECT 6.400 167.030 23.760 167.310 ;
        RECT 6.680 166.750 23.760 167.030 ;
        RECT 6.680 166.190 23.480 166.750 ;
        RECT 6.960 165.910 23.200 166.190 ;
        RECT 6.960 165.630 22.920 165.910 ;
        RECT 6.960 165.350 22.360 165.630 ;
        RECT 6.960 165.070 21.800 165.350 ;
        RECT 7.240 164.790 20.120 165.070 ;
        RECT 10.600 161.430 13.120 164.790 ;
        RECT 95.960 160.660 96.860 183.350 ;
        RECT 92.170 159.760 96.860 160.660 ;
        RECT 21.240 155.550 24.040 159.470 ;
        RECT 5.280 151.910 24.040 155.550 ;
        RECT 90.300 153.670 90.990 157.890 ;
        RECT 92.170 155.360 93.070 159.760 ;
        RECT 132.260 159.550 132.860 219.300 ;
        RECT 141.110 216.410 141.390 217.010 ;
        RECT 137.660 214.750 138.260 215.750 ;
        RECT 92.210 155.320 93.070 155.360 ;
        RECT 5.280 148.270 8.080 151.910 ;
        RECT 21.240 147.710 24.040 151.910 ;
        RECT 14.800 144.910 19.280 145.190 ;
        RECT 13.960 144.630 20.400 144.910 ;
        RECT 96.040 144.900 96.940 156.280 ;
        RECT 13.400 144.350 20.960 144.630 ;
        RECT 12.840 144.070 21.520 144.350 ;
        RECT 12.280 143.790 21.800 144.070 ;
        RECT 92.200 144.000 96.940 144.900 ;
        RECT 12.000 143.510 22.360 143.790 ;
        RECT 11.720 143.230 22.640 143.510 ;
        RECT 11.440 142.950 22.920 143.230 ;
        RECT 11.160 142.670 22.920 142.950 ;
        RECT 11.160 142.390 23.200 142.670 ;
        RECT 10.880 141.830 23.480 142.390 ;
        RECT 10.600 141.550 23.760 141.830 ;
        RECT 10.600 141.270 15.360 141.550 ;
        RECT 19.000 141.270 23.760 141.550 ;
        RECT 10.600 140.990 14.520 141.270 ;
        RECT 19.840 140.990 24.040 141.270 ;
        RECT 90.120 141.080 91.040 141.820 ;
        RECT 10.320 140.710 14.240 140.990 ;
        RECT 20.120 140.710 24.040 140.990 ;
        RECT 10.320 140.430 13.960 140.710 ;
        RECT 10.320 140.150 13.680 140.430 ;
        RECT 20.680 140.150 24.040 140.710 ;
        RECT 10.320 139.030 13.400 140.150 ;
        RECT 20.960 139.870 24.320 140.150 ;
        RECT 10.320 138.470 13.120 139.030 ;
        RECT 10.320 137.630 13.400 138.470 ;
        RECT 21.240 137.910 24.320 139.870 ;
        RECT 81.260 139.450 82.460 140.750 ;
        RECT 92.200 138.880 93.100 144.000 ;
        RECT 10.320 137.070 13.680 137.630 ;
        RECT 20.960 137.350 24.320 137.910 ;
        RECT 20.680 137.070 24.320 137.350 ;
        RECT 10.320 136.790 13.960 137.070 ;
        RECT 20.680 136.790 24.040 137.070 ;
        RECT 81.260 137.050 82.460 138.350 ;
        RECT 10.600 136.510 14.240 136.790 ;
        RECT 20.400 136.510 24.040 136.790 ;
        RECT 10.600 136.230 14.800 136.510 ;
        RECT 19.840 136.230 24.040 136.510 ;
        RECT 10.600 135.950 15.360 136.230 ;
        RECT 19.280 135.950 24.040 136.230 ;
        RECT 10.880 135.670 17.040 135.950 ;
        RECT 17.600 135.670 23.760 135.950 ;
        RECT 10.880 135.390 23.760 135.670 ;
        RECT 11.160 134.830 23.480 135.390 ;
        RECT 11.440 134.550 23.200 134.830 ;
        RECT 81.260 134.650 82.460 135.950 ;
        RECT 11.720 134.270 23.200 134.550 ;
        RECT 12.000 133.990 22.920 134.270 ;
        RECT 12.280 133.710 22.640 133.990 ;
        RECT 12.560 133.430 22.360 133.710 ;
        RECT 13.120 133.150 21.800 133.430 ;
        RECT 13.400 132.870 21.240 133.150 ;
        RECT 14.240 132.590 20.680 132.870 ;
        RECT 15.080 132.310 19.840 132.590 ;
        RECT 6.680 131.190 7.800 131.470 ;
        RECT 6.680 130.910 8.640 131.190 ;
        RECT 6.680 130.630 9.480 130.910 ;
        RECT 6.680 130.350 10.320 130.630 ;
        RECT 6.680 130.070 11.440 130.350 ;
        RECT 6.680 129.790 12.280 130.070 ;
        RECT 6.680 129.510 13.120 129.790 ;
        RECT 6.680 129.230 13.960 129.510 ;
        RECT 6.680 128.950 15.080 129.230 ;
        RECT 6.680 128.670 15.920 128.950 ;
        RECT 6.680 128.390 16.760 128.670 ;
        RECT 6.680 128.110 17.600 128.390 ;
        RECT 6.680 127.830 18.720 128.110 ;
        RECT 7.240 127.550 19.560 127.830 ;
        RECT 8.360 127.270 20.400 127.550 ;
        RECT 9.200 126.990 21.520 127.270 ;
        RECT 10.320 126.710 22.360 126.990 ;
        RECT 11.440 126.430 23.200 126.710 ;
        RECT 12.280 126.150 24.040 126.430 ;
        RECT 13.400 125.870 24.040 126.150 ;
        RECT 14.240 125.590 24.040 125.870 ;
        RECT 15.360 125.310 24.040 125.590 ;
        RECT 16.200 125.030 24.040 125.310 ;
        RECT 17.320 124.750 24.040 125.030 ;
        RECT 18.160 124.470 24.040 124.750 ;
        RECT 19.280 123.910 24.040 124.470 ;
        RECT 18.440 123.630 24.040 123.910 ;
        RECT 17.320 123.350 24.040 123.630 ;
        RECT 16.200 123.070 24.040 123.350 ;
        RECT 15.360 122.790 24.040 123.070 ;
        RECT 14.240 122.510 24.040 122.790 ;
        RECT 13.400 122.230 24.040 122.510 ;
        RECT 12.280 121.950 24.040 122.230 ;
        RECT 11.160 121.670 24.040 121.950 ;
        RECT 10.320 121.390 22.920 121.670 ;
        RECT 9.200 121.110 22.080 121.390 ;
        RECT 8.360 120.830 21.240 121.110 ;
        RECT 7.240 120.550 20.400 120.830 ;
        RECT 6.680 120.270 19.280 120.550 ;
        RECT 6.680 119.990 18.440 120.270 ;
        RECT 6.680 119.710 17.600 119.990 ;
        RECT 6.680 119.430 16.760 119.710 ;
        RECT 6.680 119.150 15.640 119.430 ;
        RECT 6.680 118.870 14.800 119.150 ;
        RECT 6.680 118.590 13.960 118.870 ;
        RECT 6.680 118.310 12.840 118.590 ;
        RECT 6.680 118.030 12.000 118.310 ;
        RECT 6.680 117.750 11.160 118.030 ;
        RECT 6.680 117.470 10.320 117.750 ;
        RECT 6.680 117.190 9.200 117.470 ;
        RECT 6.680 116.910 8.360 117.190 ;
        RECT 6.680 116.630 7.520 116.910 ;
        RECT 13.120 100.110 24.040 100.390 ;
        RECT 12.280 99.830 24.040 100.110 ;
        RECT 11.720 99.550 24.040 99.830 ;
        RECT 11.440 99.270 24.040 99.550 ;
        RECT 11.160 98.990 24.040 99.270 ;
        RECT 10.880 98.430 24.040 98.990 ;
        RECT 10.600 97.870 24.040 98.430 ;
        RECT 10.320 97.030 24.040 97.870 ;
        RECT 10.320 96.750 14.240 97.030 ;
        RECT 10.320 96.470 13.680 96.750 ;
        RECT 10.320 95.910 13.400 96.470 ;
        RECT 10.320 95.350 13.120 95.910 ;
        RECT 10.320 94.510 13.400 95.350 ;
        RECT 10.600 94.230 13.680 94.510 ;
        RECT 10.600 93.950 13.960 94.230 ;
        RECT 10.880 93.670 14.240 93.950 ;
        RECT 10.880 93.390 14.520 93.670 ;
        RECT 11.160 93.110 14.800 93.390 ;
        RECT 11.440 92.830 15.080 93.110 ;
        RECT 11.720 92.550 15.360 92.830 ;
        RECT 5.280 89.190 24.040 92.550 ;
        RECT 10.600 84.990 13.120 86.670 ;
        RECT 23.760 86.390 26.000 86.670 ;
        RECT 23.200 86.110 26.840 86.390 ;
        RECT 22.640 85.830 27.120 86.110 ;
        RECT 22.360 85.550 27.400 85.830 ;
        RECT 22.360 85.270 27.680 85.550 ;
        RECT 13.680 84.990 16.480 85.270 ;
        RECT 22.080 84.990 27.960 85.270 ;
        RECT 10.600 84.710 17.320 84.990 ;
        RECT 21.800 84.710 28.240 84.990 ;
        RECT 10.600 84.430 17.600 84.710 ;
        RECT 10.600 84.150 17.880 84.430 ;
        RECT 21.800 84.150 28.520 84.710 ;
        RECT 10.600 83.870 18.160 84.150 ;
        RECT 10.600 83.590 18.440 83.870 ;
        RECT 21.520 83.590 28.800 84.150 ;
        RECT 10.600 83.310 18.720 83.590 ;
        RECT 21.520 83.310 29.080 83.590 ;
        RECT 10.600 82.750 19.000 83.310 ;
        RECT 21.240 83.030 29.080 83.310 ;
        RECT 21.240 82.750 24.600 83.030 ;
        RECT 25.720 82.750 29.080 83.030 ;
        RECT 10.600 82.190 19.280 82.750 ;
        RECT 10.600 81.910 14.520 82.190 ;
        RECT 15.360 81.910 19.280 82.190 ;
        RECT 10.320 81.630 13.680 81.910 ;
        RECT 16.200 81.630 19.280 81.910 ;
        RECT 21.240 82.470 24.320 82.750 ;
        RECT 26.280 82.470 29.080 82.750 ;
        RECT 10.320 81.350 13.400 81.630 ;
        RECT 16.480 81.350 19.560 81.630 ;
        RECT 10.320 81.070 13.120 81.350 ;
        RECT 16.760 81.070 19.560 81.350 ;
        RECT 10.320 78.830 12.840 81.070 ;
        RECT 17.040 78.830 19.560 81.070 ;
        RECT 10.320 78.550 13.120 78.830 ;
        RECT 10.320 78.270 13.400 78.550 ;
        RECT 16.760 78.270 19.560 78.830 ;
        RECT 21.240 81.070 24.040 82.470 ;
        RECT 26.560 81.630 29.360 82.470 ;
        RECT 21.240 78.550 23.760 81.070 ;
        RECT 26.840 80.230 29.360 81.630 ;
        RECT 27.120 79.670 29.360 80.230 ;
        RECT 20.960 78.270 23.760 78.550 ;
        RECT 26.840 78.270 29.360 79.670 ;
        RECT 10.320 77.990 13.680 78.270 ;
        RECT 16.200 77.990 19.280 78.270 ;
        RECT 20.960 77.990 24.040 78.270 ;
        RECT 10.600 77.710 14.240 77.990 ;
        RECT 15.640 77.710 19.280 77.990 ;
        RECT 20.680 77.710 24.320 77.990 ;
        RECT 26.560 77.710 29.360 78.270 ;
        RECT 10.600 77.430 19.560 77.710 ;
        RECT 20.680 77.430 24.600 77.710 ;
        RECT 26.280 77.430 29.360 77.710 ;
        RECT 10.600 77.150 25.160 77.430 ;
        RECT 26.000 77.150 29.360 77.430 ;
        RECT 10.880 76.590 29.080 77.150 ;
        RECT 11.160 76.310 29.080 76.590 ;
        RECT 11.440 76.030 29.080 76.310 ;
        RECT 11.440 75.750 28.800 76.030 ;
        RECT 11.720 75.470 28.800 75.750 ;
        RECT 12.280 75.190 17.600 75.470 ;
        RECT 18.160 75.190 28.520 75.470 ;
        RECT 12.560 74.910 17.320 75.190 ;
        RECT 18.440 74.910 22.640 75.190 ;
        RECT 23.200 74.910 28.520 75.190 ;
        RECT 13.120 74.630 16.760 74.910 ;
        RECT 19.000 74.630 22.360 74.910 ;
        RECT 23.480 74.630 28.240 74.910 ;
        RECT 19.560 74.350 21.800 74.630 ;
        RECT 23.760 74.350 27.960 74.630 ;
        RECT 24.040 74.070 27.680 74.350 ;
        RECT 24.600 73.790 27.120 74.070 ;
        RECT 6.120 67.630 7.800 67.910 ;
        RECT 21.240 67.630 24.040 71.550 ;
        RECT 5.560 67.350 8.360 67.630 ;
        RECT 5.280 67.070 8.640 67.350 ;
        RECT 5.000 66.510 8.920 67.070 ;
        RECT 5.000 66.230 9.200 66.510 ;
        RECT 4.720 65.110 9.200 66.230 ;
        RECT 5.000 64.830 9.200 65.110 ;
        RECT 5.000 64.270 8.920 64.830 ;
        RECT 5.280 63.990 8.640 64.270 ;
        RECT 10.600 63.990 24.040 67.630 ;
        RECT 5.560 63.710 8.360 63.990 ;
        RECT 6.120 63.430 7.800 63.710 ;
        RECT 10.600 60.350 13.120 63.990 ;
        RECT 21.240 59.790 24.040 63.990 ;
        RECT 6.680 53.630 24.040 56.990 ;
        RECT 13.680 48.030 16.480 53.630 ;
        RECT 6.680 44.670 24.040 48.030 ;
        RECT 28.240 39.070 29.360 39.350 ;
        RECT 27.680 38.790 29.920 39.070 ;
        RECT 27.120 38.510 30.200 38.790 ;
        RECT 26.840 38.230 30.200 38.510 ;
        RECT 26.280 37.950 30.200 38.230 ;
        RECT 25.720 37.670 30.200 37.950 ;
        RECT 25.160 37.390 30.200 37.670 ;
        RECT 24.880 37.110 30.200 37.390 ;
        RECT 24.320 36.830 30.200 37.110 ;
        RECT 23.760 36.550 30.200 36.830 ;
        RECT 23.480 36.270 30.200 36.550 ;
        RECT 22.920 35.990 30.200 36.270 ;
        RECT 22.360 35.710 30.200 35.990 ;
        RECT 21.800 35.430 30.200 35.710 ;
        RECT 21.520 35.150 30.200 35.430 ;
        RECT 20.960 34.870 26.840 35.150 ;
        RECT 20.400 34.590 26.560 34.870 ;
        RECT 19.840 34.310 26.000 34.590 ;
        RECT 19.560 34.030 25.440 34.310 ;
        RECT 19.000 33.750 24.880 34.030 ;
        RECT 18.440 33.470 24.600 33.750 ;
        RECT 17.880 33.190 24.040 33.470 ;
        RECT 17.600 32.910 23.480 33.190 ;
        RECT 17.040 32.630 23.200 32.910 ;
        RECT 16.480 32.350 22.640 32.630 ;
        RECT 16.200 32.070 22.080 32.350 ;
        RECT 15.640 31.790 21.520 32.070 ;
        RECT 15.080 31.510 21.240 31.790 ;
        RECT 14.520 31.230 20.680 31.510 ;
        RECT 14.240 30.950 20.120 31.230 ;
        RECT 13.680 30.670 19.560 30.950 ;
        RECT 13.120 30.390 19.280 30.670 ;
        RECT 12.560 30.110 18.720 30.390 ;
        RECT 12.280 29.830 18.160 30.110 ;
        RECT 11.720 29.550 17.600 29.830 ;
        RECT 11.160 29.270 17.320 29.550 ;
        RECT 10.600 28.990 16.760 29.270 ;
        RECT 10.320 28.710 16.200 28.990 ;
        RECT 9.760 28.430 15.920 28.710 ;
        RECT 9.200 28.150 15.360 28.430 ;
        RECT 8.920 27.870 14.800 28.150 ;
        RECT 8.360 27.590 14.240 27.870 ;
        RECT 7.800 27.310 13.960 27.590 ;
        RECT 7.240 27.030 13.400 27.310 ;
        RECT 6.960 26.750 12.840 27.030 ;
        RECT 6.400 26.470 12.280 26.750 ;
        RECT 5.840 26.190 12.000 26.470 ;
        RECT 5.280 25.910 11.440 26.190 ;
        RECT 5.000 25.630 10.880 25.910 ;
        RECT 15.360 25.630 15.920 25.910 ;
        RECT 4.440 25.350 10.320 25.630 ;
        RECT 15.360 25.350 16.760 25.630 ;
        RECT 3.880 25.070 10.040 25.350 ;
        RECT 15.640 25.070 17.880 25.350 ;
        RECT 3.320 24.790 9.480 25.070 ;
        RECT 15.640 24.790 19.000 25.070 ;
        RECT 3.040 24.510 8.920 24.790 ;
        RECT 15.920 24.510 19.840 24.790 ;
        RECT 22.920 24.510 23.480 24.790 ;
        RECT 2.480 24.230 8.640 24.510 ;
        RECT 10.320 24.230 11.160 24.510 ;
        RECT 15.920 24.230 20.960 24.510 ;
        RECT 23.200 24.230 24.040 24.510 ;
        RECT 1.920 23.950 8.080 24.230 ;
        RECT 10.320 23.950 11.720 24.230 ;
        RECT 16.200 23.950 21.800 24.230 ;
        RECT 23.200 23.950 24.320 24.230 ;
        RECT 1.640 23.670 7.520 23.950 ;
        RECT 10.320 23.670 12.560 23.950 ;
        RECT 16.200 23.670 22.920 23.950 ;
        RECT 23.480 23.670 24.880 23.950 ;
        RECT 1.360 23.390 6.960 23.670 ;
        RECT 10.320 23.390 13.120 23.670 ;
        RECT 16.480 23.390 25.160 23.670 ;
        RECT 1.360 23.110 6.680 23.390 ;
        RECT 10.320 23.110 13.960 23.390 ;
        RECT 16.480 23.110 25.720 23.390 ;
        RECT 1.360 22.830 6.120 23.110 ;
        RECT 10.320 22.830 14.800 23.110 ;
        RECT 16.760 22.830 26.000 23.110 ;
        RECT 1.360 22.550 5.840 22.830 ;
        RECT 10.320 22.550 15.360 22.830 ;
        RECT 16.760 22.550 18.440 22.830 ;
        RECT 19.280 22.550 26.560 22.830 ;
        RECT 1.360 22.270 6.400 22.550 ;
        RECT 10.320 22.270 16.200 22.550 ;
        RECT 17.040 22.270 18.720 22.550 ;
        RECT 20.680 22.270 26.840 22.550 ;
        RECT 1.360 21.990 6.680 22.270 ;
        RECT 1.360 21.710 7.240 21.990 ;
        RECT 10.320 21.710 18.720 22.270 ;
        RECT 22.360 21.990 27.120 22.270 ;
        RECT 22.920 21.710 26.840 21.990 ;
        RECT 1.640 21.430 7.800 21.710 ;
        RECT 2.200 21.150 8.080 21.430 ;
        RECT 10.320 21.150 19.000 21.710 ;
        RECT 22.640 21.430 25.440 21.710 ;
        RECT 22.360 21.150 24.040 21.430 ;
        RECT 2.760 20.870 8.640 21.150 ;
        RECT 11.440 20.870 19.280 21.150 ;
        RECT 22.360 20.870 22.920 21.150 ;
        RECT 3.040 20.590 9.200 20.870 ;
        RECT 12.280 20.590 19.280 20.870 ;
        RECT 3.600 20.310 9.760 20.590 ;
        RECT 13.400 20.310 19.560 20.590 ;
        RECT 4.160 20.030 10.040 20.310 ;
        RECT 14.240 20.030 19.560 20.310 ;
        RECT 4.720 19.750 10.600 20.030 ;
        RECT 15.360 19.750 19.840 20.030 ;
        RECT 5.000 19.470 11.160 19.750 ;
        RECT 16.480 19.470 19.840 19.750 ;
        RECT 5.560 19.190 11.720 19.470 ;
        RECT 17.320 19.190 20.120 19.470 ;
        RECT 6.120 18.910 12.000 19.190 ;
        RECT 18.440 18.910 20.120 19.190 ;
        RECT 6.680 18.630 12.560 18.910 ;
        RECT 19.560 18.630 20.120 18.910 ;
        RECT 6.960 18.350 13.120 18.630 ;
        RECT 7.520 18.070 13.680 18.350 ;
        RECT 8.080 17.790 13.960 18.070 ;
        RECT 8.360 17.510 14.520 17.790 ;
        RECT 8.920 17.230 15.080 17.510 ;
        RECT 9.480 16.950 15.360 17.230 ;
        RECT 10.040 16.670 15.920 16.950 ;
        RECT 10.320 16.390 16.480 16.670 ;
        RECT 10.880 16.110 17.040 16.390 ;
        RECT 11.440 15.830 17.320 16.110 ;
        RECT 12.000 15.550 17.880 15.830 ;
        RECT 12.280 15.270 18.440 15.550 ;
        RECT 12.840 14.990 19.000 15.270 ;
        RECT 13.400 14.710 19.280 14.990 ;
        RECT 13.960 14.430 19.840 14.710 ;
        RECT 14.240 14.150 20.400 14.430 ;
        RECT 14.800 13.870 20.960 14.150 ;
        RECT 15.360 13.590 21.240 13.870 ;
        RECT 15.640 13.310 21.800 13.590 ;
        RECT 16.200 13.030 22.360 13.310 ;
        RECT 16.760 12.750 22.640 13.030 ;
        RECT 17.320 12.470 23.200 12.750 ;
        RECT 17.600 12.190 23.760 12.470 ;
        RECT 18.160 11.910 24.320 12.190 ;
        RECT 18.720 11.630 24.600 11.910 ;
        RECT 19.280 11.350 25.160 11.630 ;
        RECT 19.560 11.070 25.720 11.350 ;
        RECT 20.120 10.790 26.280 11.070 ;
        RECT 20.680 10.510 26.560 10.790 ;
        RECT 21.240 10.230 27.120 10.510 ;
        RECT 27.400 10.230 30.200 35.150 ;
        RECT 141.620 20.710 142.580 21.400 ;
        RECT 141.710 11.180 142.050 12.010 ;
        RECT 21.520 9.950 30.200 10.230 ;
        RECT 22.080 9.670 30.200 9.950 ;
        RECT 22.640 9.390 30.200 9.670 ;
        RECT 22.920 9.110 30.200 9.390 ;
        RECT 23.480 8.830 30.200 9.110 ;
        RECT 24.040 8.550 30.200 8.830 ;
        RECT 24.600 8.270 30.200 8.550 ;
        RECT 24.880 7.990 30.200 8.270 ;
        RECT 25.440 7.710 30.200 7.990 ;
        RECT 26.000 7.430 30.200 7.710 ;
        RECT 26.560 7.150 30.200 7.430 ;
        RECT 26.840 6.870 30.200 7.150 ;
        RECT 27.400 6.590 30.200 6.870 ;
        RECT 27.960 6.310 29.640 6.590 ;
        RECT 33.860 5.700 34.460 5.750 ;
        RECT 101.380 5.700 101.800 5.710 ;
        RECT 33.860 5.100 101.830 5.700 ;
        RECT 33.860 5.050 34.460 5.100 ;
      LAYER met3 ;
        RECT 128.060 224.685 128.660 225.235 ;
        RECT 129.810 222.500 131.410 223.500 ;
        RECT 123.810 219.275 124.510 219.925 ;
        RECT 92.160 217.500 127.560 218.400 ;
        RECT 129.860 218.000 131.360 222.500 ;
        RECT 90.230 208.875 91.020 213.045 ;
        RECT 92.160 211.395 93.060 217.500 ;
        RECT 126.660 217.200 127.560 217.500 ;
        RECT 126.520 217.000 128.110 217.200 ;
        RECT 126.520 216.985 141.430 217.000 ;
        RECT 126.520 216.435 141.440 216.985 ;
        RECT 126.520 216.400 141.430 216.435 ;
        RECT 126.520 216.300 128.110 216.400 ;
        RECT 126.660 216.230 127.560 216.300 ;
        RECT 92.160 210.495 93.110 211.395 ;
        RECT 95.910 210.575 96.910 211.525 ;
        RECT 92.160 210.440 93.060 210.495 ;
        RECT 97.860 189.500 124.355 215.500 ;
        RECT 137.610 214.775 138.310 215.725 ;
        RECT 90.230 180.755 91.020 184.925 ;
        RECT 95.910 182.375 96.910 183.325 ;
        RECT 97.760 162.300 124.255 188.300 ;
        RECT 137.660 187.200 138.260 214.775 ;
        RECT 124.710 186.600 138.260 187.200 ;
        RECT 90.250 153.695 91.040 157.865 ;
        RECT 96.120 155.455 96.900 156.235 ;
        RECT 48.560 119.700 80.055 145.700 ;
        RECT 90.070 141.105 91.090 141.795 ;
        RECT 81.260 140.725 82.460 141.000 ;
        RECT 81.210 139.475 82.510 140.725 ;
        RECT 81.260 138.325 82.460 139.475 ;
        RECT 81.210 137.075 82.510 138.325 ;
        RECT 81.260 135.925 82.460 137.075 ;
        RECT 81.210 134.675 82.510 135.925 ;
        RECT 97.760 135.000 124.255 161.000 ;
        RECT 132.210 160.200 132.910 160.225 ;
        RECT 124.710 159.600 132.910 160.200 ;
        RECT 132.210 159.575 132.910 159.600 ;
        RECT 81.260 24.970 82.460 134.675 ;
        RECT 81.260 23.770 142.690 24.970 ;
        RECT 141.490 20.630 142.690 23.770 ;
        RECT 141.660 11.205 142.100 11.985 ;
        RECT 33.810 5.075 34.510 5.725 ;
      LAYER met4 ;
        RECT 128.105 224.760 128.190 225.215 ;
        RECT 128.490 224.760 128.615 225.215 ;
        RECT 15.030 223.500 15.330 224.760 ;
        RECT 17.790 223.500 18.090 224.760 ;
        RECT 20.550 223.500 20.850 224.760 ;
        RECT 23.310 223.500 23.610 224.760 ;
        RECT 26.070 223.500 26.370 224.760 ;
        RECT 28.830 223.500 29.130 224.760 ;
        RECT 31.590 223.500 31.890 224.760 ;
        RECT 34.350 223.500 34.650 224.760 ;
        RECT 37.110 223.500 37.410 224.760 ;
        RECT 39.870 223.500 40.170 224.760 ;
        RECT 42.630 223.500 42.930 224.760 ;
        RECT 45.390 223.500 45.690 224.760 ;
        RECT 48.150 223.500 48.450 224.760 ;
        RECT 50.910 223.500 51.210 224.760 ;
        RECT 53.670 223.500 53.970 224.760 ;
        RECT 56.430 223.500 56.730 224.760 ;
        RECT 59.190 223.500 59.490 224.760 ;
        RECT 61.950 223.500 62.250 224.760 ;
        RECT 64.710 223.500 65.010 224.760 ;
        RECT 67.470 223.500 67.770 224.760 ;
        RECT 70.230 223.500 70.530 224.760 ;
        RECT 72.990 223.500 73.290 224.760 ;
        RECT 75.750 223.500 76.050 224.760 ;
        RECT 78.510 223.500 78.810 224.760 ;
        RECT 128.105 224.705 128.615 224.760 ;
        RECT 129.855 223.500 131.365 223.505 ;
        RECT 14.990 222.500 131.365 223.500 ;
        RECT 33.360 220.760 34.860 222.500 ;
        RECT 49.255 139.200 78.865 145.005 ;
        RECT 79.555 141.000 80.035 145.640 ;
        RECT 90.090 141.080 91.090 222.500 ;
        RECT 129.855 222.495 131.365 222.500 ;
        RECT 123.855 219.295 124.465 219.905 ;
        RECT 123.860 215.440 124.460 219.295 ;
        RECT 126.555 216.295 126.560 217.205 ;
        RECT 128.060 216.295 128.065 217.205 ;
        RECT 123.855 215.100 124.460 215.440 ;
        RECT 95.955 211.500 96.865 211.505 ;
        RECT 98.555 211.500 123.165 214.805 ;
        RECT 95.955 210.600 123.165 211.500 ;
        RECT 95.955 210.595 96.865 210.600 ;
        RECT 98.555 190.195 123.165 210.600 ;
        RECT 123.855 189.560 124.335 215.100 ;
        RECT 123.755 188.100 124.235 188.240 ;
        RECT 95.955 183.300 96.865 183.305 ;
        RECT 98.455 183.300 123.065 187.605 ;
        RECT 95.955 182.400 123.065 183.300 ;
        RECT 95.955 182.395 96.865 182.400 ;
        RECT 98.455 162.995 123.065 182.400 ;
        RECT 123.755 186.000 125.960 188.100 ;
        RECT 123.755 162.360 124.235 186.000 ;
        RECT 123.755 160.800 124.235 160.940 ;
        RECT 98.455 156.300 123.065 160.305 ;
        RECT 96.120 155.400 123.065 156.300 ;
        RECT 34.860 128.400 78.865 139.200 ;
        RECT 79.460 140.705 82.460 141.000 ;
        RECT 79.460 139.495 82.465 140.705 ;
        RECT 79.460 138.305 82.460 139.495 ;
        RECT 79.460 137.095 82.465 138.305 ;
        RECT 79.460 135.905 82.460 137.095 ;
        RECT 79.460 134.695 82.465 135.905 ;
        RECT 98.455 135.695 123.065 155.400 ;
        RECT 123.755 159.000 125.960 160.800 ;
        RECT 123.755 135.060 124.235 159.000 ;
        RECT 79.460 134.400 82.460 134.695 ;
        RECT 49.255 120.395 78.865 128.400 ;
        RECT 79.555 119.760 80.035 134.400 ;
        RECT 140.770 11.140 142.130 12.040 ;
        RECT 140.770 3.900 141.670 11.140 ;
        RECT 136.170 3.000 141.670 3.900 ;
        RECT 136.170 1.000 137.070 3.000 ;
  END
END tt_um_urish_charge_pump
END LIBRARY

